`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
N9UGgKGWxj0dC5CZbJU17jocbWLNhNOTb3aPljvAtUlt1z70r0bgwKQFhJ0YenCTxVkTnqKOkuGN
0HZ2B5qrUQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FmEHqkkbGHYGnl8i3ASmJSbcE71EsvvIpV5j21oFdm76AMUN5Mrzc48nnQgtTmansEs60PdK3xP3
QToOegG1CtWssFGK4djltTWGP8CMTuVs1sQZIbRiIgP4zCKykzPHw7awLfmdNAvyT7c9P4/PxToV
7s7CTIYrcwEuF/mVIgU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JkcK+z0zcFSMCI3qblNs01iANwT/eBRnX8RrMwhUtfXOWjmJt1ylkizXaOcASnqi1PbASAdPaDgw
P1J9CF1xBro3dKkiZjDq5gLqLdCNMq+Qhoa9QaLLhY9nftxquC7LiM+S/DXIUdSrcb0Ok5jDOmfP
V9i6hz69i26VdK1rRRZ6Ufc+YKCO3+9CH/DU1mMgy3zQmxaTQI7sRCM+dTMwgVeJ+eFXieGMI6Xf
OPNeuiLXFepchWpFvkzMmto0Lr4oFXtQOtqSosIlSpHh7aJ9/J++OJwXD668nRMsaoNAvdjaf4J8
+zkQI7domt4j02cvx1P7c+bAvgxT0khT/5b4pw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CXzYa3CwhfcjP6YB70R+BJ8KOoGZ77fl+2VswrlXcD5x43kUvWe/ElpepDS4x2qEygwPbO91SI/g
qOY+YkHj92X5e7U2EqsIZpC1e5G289b5dr/uGJCXwEHWECmWBV4DXlUUSSKb8ONEl4beLI6Fqp5l
DHVXJsJLI5jQjG5HxgI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rr1CKBq86wNPNUMynPvJ74u4cIprzV+nHUFd8Q+D1/lqbRYit3k4lb09yQrk1//8dSAeItZtjDHN
8NpKAmf6GrwUgcOwDoiFv5ygl0sxoFhSFSjmZ5d+FTVMo03Ap8x+qIIfb/qu4yqJmyi+o5BWnhjw
y7lUkCpB5xY4vOKIEO4VBXHLqnjkeNnBn16tp7EyT2EvYVuWG/NXk2enSxCxirrsTbqC8aXzU1qP
k8etpOb8byva5iJS2rujLsGm74TsBqGbYeyU7oa/Sp1tOoA++dBl0LZj68LZL0vWSHbOUvDCUhhZ
4kf5A0WrlrbCE/P2Bf9lhWp2nD973ZtMWeIkUQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vefzraaMaUcgUXELf03iKU/IrUYEauhHMQ2CqLgU8RXKO0BanYiY2ubtLEx6pUdzYU7VnKC4/T7N
y/25gTbiM8zets9B4DhtG5ZVGYrZOvVCHivzcp6tAPjnvpGV5ato037yPaZIv9tS6tjPiOVM6tvZ
G5FHuRav0yX2SDsSmpUXBalAzIH5YLMyDNeENoO7N8Ujj6SyiMUSY18VQKBNXl+mU59c9imzZrLS
hwtL7l17GDQE/uLsXgEnJmp8eOEBrNvR5/mJhInflqCG9740hURij7gOm4ofuKxI05r2kiqQJUZ8
tZKvIg9X9RGMPZFmEiPZmo8beZ6MQDhKwmx0QQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16928)
`protect data_block
G2IN9yVKGesaBlUHEkdk5UwqOJU5RHaVc9xmjq8Io1plLU5HToNTA9RYnc1v91VRk0SEgluCs1Ik
XN47yiJRRH+B4fLX2JBlE1fMNlz+GlTmqV9+5UW+lQkF6KvIkmM4ZjPx46UlM7hRpvfH4RgVBuFT
Iej8zS7PHDr/bTRbQH6gd28+w96Im82fZ/lncfcf16rmwOPXOaxxYSZBVcOLp9lOf2eS713SS2MR
cnhbhv/vpPEy8tV7DyriTeOI/OKZsBEt7wrFHQgn5zRfnopA3k73asTTHJF1NKDdckxC/VvrChJq
cZdy63JikvXWO38qar1sQluq0+DIWJcGVIrUNwtn+MQcSDyDnrNgjSo+WkqXwRylj2uu/Uak3h3y
aTDqeu6uB1vUiATsjmz/tNj0IDNaxQcx6m9nwaGc4fH0o+nMasNtxCi5r4D8REBXtmu4fqtG4sdX
oS/OUSWZUu5idoqYO2pmF62N1YWEZ+U8Y2WBVcYj7otMKLxif2Av+K3ZUFR3xd8HtdBRhqP437Rw
xt6s09eOoQ3tcE9f/Em3FVIQsSuVUCM67qERv8adFUb5lh/NlkR8iW4hrvjgVqgcIh7kowtUsiyY
zekgqpq/YezBfqC/U4vB74OJ7AXi5HwZDkBwaeG09rBUPJAYHVQVRusToFsiJHWV2QPBUbNhbutO
zne4FczQclMdtLKW0VHOWrm+0WSIFkRunhgQECjeyqJjVzUqqnF3qtujbcSOh2bPLep1BcemK77t
/dseFr3c/nADmTLh6oZODxPjIerpS9VEYWVP0m+Kcxn3nWHdq71DJ3R95Oh5IoZx1jjLHsXvq5fL
Xsh915XULbSLJJbtKsiLxFfyldN3ghoROY5SH0XftBOqan0uK4PiGWWe54QgxekwqQuqLRrle6SY
NOS/NOE7vMrZuRLl0K+MtBLUl2x17PDwJprb2RoQN9aXA2KkP8dqIiMR7hX+TzvPwB43yB1OeWZ7
hkcPTcDYStdhgp8/VZd3Z+VXvBw9vXJXeiHujuh2uTKfTS8t/j1f0FqXKTUG9rOMFDMoFcOgB/H7
eXnvaLKrpTbTGPTuOu1qqezsprEtQED1m0uGE3m6jyDs7RWK83s0q5vhzOxWSgEvP7t/oA/SCcCR
gmUj1SVZHowIJif7cCRy2LNRIixYv+jeCLysMo0TK4eijkaxYiI0RFkOXhsHAIJ2kzGDcLH4NPqm
w8nHjGmrU6LYAdkcqDkUqvVuwBEJv5PdKNlhwP6q5B/VXafPBCL2c9wiVaORSSb4Un/tIE9whLav
2Kmk0n9ThnbIVGGNYATYfxfhnIeSMpIZZZZ1xk5T1suCCHkqstM9FDjwW4+i56GTymmrcwZ+B0bL
qv2/34WaOAyu7cLX5HgzYMr2VZz7YEhgAx9KirvzlgC3Ab0MDTylF3XpPF+Sjqe/yh/rzWZ9D63L
R9fhem6Ehvv2+t83LzOVx8zxeWqMHBrm7ZIruYBbHCRPjgqffK6tACpTxV8fy8irN8r5NGURIgJW
eCPxUOhAMTvtZmO5J7ugW9UUxew6xS5fziT/KySjWP14VsYAq680BN1fRPCqRPVn4hcwupzylQTA
0KMC121RjHwlYIjMstNOBscemZBTvJNgvpEGJ1S1COIByajHq0VdQlgYEbLen8ZbaTAGLINmBjXB
iM/A5AdGf5j3WrU+UjLLvElT2MCpl4/S6hwS/2WBlWsF3aArqtvgmEDyFEE0BtxADFs7Hu8P9Wir
1JVr5sOouG5Ba2eUb9FtfIigdFj3GekAfj+nX+JMPpRJKYuC7i81V6cqTyHDArHdAbXeDhAltbyu
YB8+KGcklLf2Krnyzmq0AxUztm5yzL6zcSmGtGF3kRdOLELU3VadmAnF/MJvDz5OKR57oirgIuuP
9D99zRx74xD7OhG9wgUF+3nd1b5OI3llGEuRkBmtEJrnAUs5mzS4T60RX4iBRE5Kb1QBJUjltVQh
XD3uh2vYy0WxJS1zj99d/crFPADizCHvVVdFmgyaqMmeKHZ3MZrfjdL165CPJtsrRZHwFDCJUQUZ
AucHcheITHh14qxvkbGEqo9E29Y3B1fzLTf0tFiS2I2QDBP5Q2Usk5D87k9B8cSW81L4JV0lAqdB
MIHD9kJGxyE3LHjgtiZr7oSXe7E3a3SQaAGxz5zsZnAtyZqIvx8Zdy1k/bC7NuN8qkE6MDwyDqAm
IP3h2ooqwAwLkaDTvdVSg2TsdDO0Btt+OU0WwWiEZMvc0Uc2XNIEjYfOasvmqjvGD9sevx9c4fyk
aMaCKxmqO1V87r/28+Pl4DdLPNWOUNQJWVr03G4VvYdPT6r2LYGAmno47SboPCEPQGX8v/LSgRy2
XLLBILPg/25Q5cZBw84VgjFEZPqB8Wr6ioFBQUJo7U4v+SEwfODPNl2E6XaEQRyEyC6URyg6DTlc
9FebK7rVtPwjLAap9b1TpWb2StqQI3sxorqxcxN7gL0u1JpF52IG0k9oK6MrIjpR8Ot4mdbFwkCe
75aR6XGff6xItSqzaWL0fDb00DJEFEl3obBQ2cRshqo3MjMCLkt+J2yZlFonazK1KLwj28EbZQW6
CcCmjX4HxBXUeUBDvspnUVm2yBim12IQ2QbdelBrdhgUKNnNXLsEBqco+wjK/ZZ1MaGCnH6WeOs0
fWITNplYtyEkg6LUV+tZt5dWW+vcfWY46BpoZju2GKT0+YxjTT3ADCrBGURXP9WQwuNGm1yl8Ron
j6Zup5zUqV/ceHTvEwpPVYUEP3YsHYiG/oK61jz9kbR8s4A4IYh+7+4WYV772fHBCCR6qQ1PExzY
c1h/TeqhwmzcGup7Wgp3E048OfKSxd593qdNkIItjdKRHaaHHjeXs9IHaTOQhME7MiMwwDZAnhyd
TGu2Iy3YV6ZJ/oM8f653hYIcfN78S5rvUBDhtNR3kwROaxgPnolEn56peX/86dapZsLGeClnVKla
bQyNkZDg2VNMK5o6lTl7fODnK04St4uIkE58VnWcV9E62cqgjfT/a/mII9RpYhe6n8xZ/SQHemnl
JK0OjR42ohhRMNGf7sr+Fb7fyH/E7mvDp60UQLUnQRMUiaoxUB2coPD4k9qr741g0807AtH5APwZ
SqbGSe7InRwGCcYs6pn7mZWTyyeaCwI+f250ZkLyb5ZlEjmE+qF/n3+hGnoTt/S7vD6dozZmHmz9
h/vHc/ql+PPAEH8cLiODE29cGvkd5/9dRrAdkIycVUaHW5yM4drCw3SH2rjJLeguHWDZEwguVlqn
UjoFjvsJSXbj897mP30BruQDarWrPBIZ8C38G5Hc4jiy9DbCh21CStgOjJmYnxA+3H/JJizGozc9
0e/eIDhdZy+mLZ55ntYUaTEg5MlXCwIJXMD2xpr4T1HrqN29couCaOek83ox5QWdTFZkkZnslyXa
3AcwjuRJOyPGzSe9GKILel23hM7P7KbbMzZQjvtz3m3pBS2auET5tLJznHb9S01BQl/ScqeC4bmA
kSoJkHa3Usv2d2MNnsZIhkDMh4yPvJgRa02RlqMQ5ZmpfpG3nQImONoVLeCs9ljWIaovJIS9KbNJ
Kmx8BLdeQmccSfXbZdABPkJPqkWf5qeL62m6Q9VUi7THqEKMef9rZ+u28hKH6jzCbKPKPRh+TDCW
X5LVqGD8Nr2JBQaA8kSPtYov+Eb2HJNhpt8orVKjKQX0X/jsb7hdlfsP3Hvv2WMLnIiUATtF7X07
w3OyLXryTCQqC0FQ4uEeOA465zDWo/Gd5yxsY8XEGxSJcz/or1z1Q1HT8ZVIH/QQ3gHNsABDF99c
a3N0vEHUPWJN4uRXrSetU1bAyUUHjj5+Dx3oTexSqvpCRa5xkQdS1mPZbCsphqH+/V/R7eTFNA16
IhzsyVfMwE//pljBHe4446kl9vXHEN+LuXY5tiodeHmSClQYmnB/rOgejhyCct3Qkr5kRJ40QO4w
AO3ONneEbAZI0JwGVki5iqV+OiRUUYJYQ15UjQ8J4BCNvTebuqSjWKXfF5NWYmbyYxYuEU6GClZh
LB8CcM+Lr9oLz9VCVGYcHY6c15uTCRXhpwsCvKCp52lgAv+WMOhwAXA/AfvrSeiISWt6mrEWNp/G
sQOhZaT4Ft7Snc2u0nHfobFRuGj9djUrxOsl6U88Idv/2XGn9Rk4DybKxWcTkJqpNWHOhIg66JeQ
fm4DDKwD/GsrPapUh4Yez3UXxDMM4PSBgw2lVNmicvjvX8w/L063D9n6ETX3EgqrIYRCWaokfpC/
5sPRZX7GHljYDk5g6G9qC5mWvs9Vs7PN+dl0iYGHYaDRLvqjggoV2Ftlz98x+8r7MGkO0J7vNpU6
Q+T3dl29KjHL1YJwXPICflQ4gfg7Nd1ezVAS9nPkupeZeR53j8KTY//3W0AOq/11/bajyVitrh2H
ozJxqpI0mqoYwIprkCBGMkk5zYuuC+fKzkSlZ3mr5pLdbAxJgYnEOZZiLTkvLtzd0WDqCeQON+We
b6xO61QSUaILK5UwQS5cTmTZRValfaeFo5lMqgSGKXdcJvLOC451AfOf6KxTx0oEyL30rbrpQ02+
fEE8e3tQmrlfpIxcZqRu7Q85sk5EV6CMo78EkvvjS6ORB46S/547OiFJALFcKdOAJD2+UyQ9qnYe
XKgQVxiGyOrgjsofgbaTePkPfysKycqaUZpiEcu88rrXst9B23GGsnX9BJMvhJiuX2FcPQBh5x3v
/2no/t92GxL2v6jC6RsBn7/2PDWeYSgej4tkjOjD2vki61WDtE37DUZSNLZgEOr/cFegguOzTWnf
piHa6SA/eUNBbmk/UoxrZKZZpnKBCazv1ibv3A+VA11ZtSDd3vPXvL3jy8U9nAHAwI41G2ykYBvS
PRgsnU1fKr0zjRKxoWK++ca29pX6nzCtUkE0O+QCwLuoC7HtzRHK30uhvd4yW3VNQEfwannYC0hj
jNZXea606024UCVAnzO0YE0l+oZRVFeMWmJXY0DRsgXV4+ji90hVHeigv43aAqotnOi2syFWnf/J
/w74tlBscesZrNlPVf1QtE1esl/UwyLG5zP26atzaiPHeAVkSUtNIhKmfOJjnhed3X+o+fpOYRls
FQTIrxTAjmu0LFZnpbidjDsA2TJPfPCBRZ+LBOJNTuO2E8HsVjAF9RqxDsLYefdkD7KXAMHFN4NA
1cywK2hTdG2OfP7tcGIHHv0HlytS614j3TesPzM9a6Uqyhh71fSxYwUvbMAacgn68InfmHRrBKr6
guNWQQjrz/qNB9ZOG5uWZnLAbozT0f1iQX7CqskXjfUodh5pOGXKJtdDlBHHMz61QVJhtyaVXDNJ
zO+A/2GQV27TwFhbE97SM9pBC51/x4yKb0ky4xa8KSfkQkcPgOl1AI+cQjFnAuKw85UIPtEvMl1j
4cZyRFSV2BYKaqpyR0JX+92gaw3oV/0rYY0nb+YQpN6WzlRVY0237ei83LGq0JsLC9iy96ABtU7R
xoqyHqehzbpm4JmpvEV/yo0xAdJuUaFlNmBmGTBDrRtpw4q+zFv/ph4AVPdiS3z9/RtRx4gVQ3fz
YCiLTHEbU99HCEZD+ok5FaIHrHO4VpDdcLzrZpJTi/6Z+R5jSZ4upyyT98ZUQKig7c3oCVDhwNQQ
71fo84biPLJLXjgfeO9GAxXLT/utE6HYApHr5YeOlRpi+Ox3t6MVmO9yD9b41w0MC+4YAaRGXWGd
ORJiJsWeRuizl6uu46Ie5v8jKo/wtndT5VOYWIdyhdPygO6uaNO5G/Sc3H6BvMvJ2kzEachXihNW
3pB2DEdxXZasmh70/Vnz+K6uJqd2HPUfGo8RG74UK8sY2Nst1zH8UnT/J0anJ9/WRvi/yw8imEun
ucUJLxA7IKCM/8rVhX2z7MZsHwrHsW4mYDiusb+LusnY8DVabF6XcNirD3keuwxOL7UkqinXc1rw
N6vc3G6rguFX7ELitl8WWH8Fneu26U5uHddH7gTbTRS+y0yqv+dH2iJHrbRhTiEaq+Hp2eddUERF
J6eKBaCoO1yGMoa0bkp09wlOGAFIIQRiEOiQtAxsTT/Ywf2EJcOD7JjUcY9R3Lpx3jpqhR4iEf78
uamJv243aNDMsVGr0sVNrOsLf3IG2RqlgJM3XxIG0EVv2xntlfTNaYozXqFEsd+v8KbLa8jyEkM8
ILNbFEyvkhdTZ4Av75YftAOGb+blEAuqweHiMuloZa2fM5pCuZuiqQLDq/N1Q7E/j7BCHAXjejhA
VqTZcKGTijWcHC+UDuBgsuuy3MHER/uTyYmuwEzSEYI1OMlmYQeA7LhkHwkswOnMJdA5FNS352pP
bqFheBzIHXdBw4rFQVvTdFjHTBx60cFRpOlUUu5JlBatF30j+XuN58MLzsQANjHLdXlui1CPEKMg
NimWZ1X6UxxzhB3KZMVOBZ5D/oXjFRzl5lT/pGomrox+Yz36N3Qv+1hhNMLUeeQGYRWdwsMsDl8R
pSBFh+vphkRgoGE1EGFWXdwRJYZqYKpkC7BIE1bso6ud36ue8XtreCr9YacfucBzcHOkpZkmkZs+
0oI2ZDqQqkgcQsfTjIAxZRUqj8AjtsKWoGYZcwnRWKbMi7b7lGXfER2vAPFDJvnUd5IWNKn9O7W6
OIKESZFlcGeklcS5dq69rcO12CH+NfW33xTlo5exYgzIvesMsyz8mFT6uJPaebrK8zg76uhpo7Uj
GPqDuAR65ZrrKLzZGwmkA8Ux1MT/nRzQNsaJQ0X0TExsp6AhHIJ15SGyTIbyrqNcWrJ5i8GHUd/9
soSJCI2ElEaPMPBLlu9ijJ7HBLxdaBE5XJkhx7qefiBts+yapg6pQf67SQlCP7Upagp3HDX3XNYi
iTmdnDW/ds4qWgrXAsb6NdRAXUll0ewl686u+K5i0e9Dta9RAgEzY9HplL+XiN8lAJ8UwW+MrNna
0QU7sMZr/H5h/v42mI2CGLw3X/3APONfj13V4pNbrxQ6CRTwypAbhFkbgv9Ch7M5eDMx7chtpqe+
73aRmiF0wp46yjKwW7VdSmiRLpaHclBi9pg22l0NJ26OF2QwTLXU4Bqog265MlPSVqX7TzJ5MpF/
34PiXhTtt1rJ+jwaBiZEZMXLtSVLOJwEbXvu+dwTmncnROvYKuXmc6JaacT3N9grlGEU9dWplE0Z
y8E6zNcVNf8vmEeWjIkrJrtt9VzgYkCSRClGPawszB+fLhWWohefhQ4cWwBKmpFOehlEFVU3MgeX
ymjDXuKmgsS1XkxI+t/kaQaZkpbhzYE2QV0gXURUIu0O/V+ziNkAtYZ8BarlCMh9mSl6qgiOePxW
o4BTJF98BicTeTMcCM7RfSEcLFIwQypY/mt4gsYbNf3RWcqbtMNNzA7kpSGC73pXvfmS8HfuAiDf
xTMUVxOHw+rUFlY63fJ8BgctTzqOyOrze84UFX6VEgLbBqzxHkVedHAWRh+VRyc1YvT6F7KS7SR0
4mZJ8BhdMbkypz73NLQxDCfir8uFnIswDZX8/V8vrvyQq1mu5NPMSZ7sQXNaG+C9/AfKiNJAaVAd
pg8T6AG6ZV9R7muCtY6YrUYKvTQDIoIq8crvi9lMnAPsS9IYcRNEkqeMLeogdI7w0JnP9ifrGS/b
zun5edmtOSz3m9N7ekrG6++vesSTHettgAxSSAvvhXVAR48Tmg3m6+hrsjsbSXwbjOIUvWsARFzF
Hqtf1y9SlIGfQrKgQ6OMgt/rb9fBr0E8OxaXkTZuDbQrKDclDVZiLMFtbGU42B3Hjsk7Hqs/ieo1
KqZN1dJIW1tmkC0aVY74d9HwFe7pF9b/4S+r8onEcfqhlGap72goh1RakBYAp5m4vL2xaIjTg5hm
ZyY/j4rsxunzsTZtd47NDmKLQ6Qkf/Tt0NCdR1sSc9jXkqhQIQef9khyspCGiZry0um1pX08J++x
tULr9LqzPvZvq1+KFc+RKiuHG5W/Prgqdg4n7+jsvG9w6d3alcdWOTGLCDoRxH/JtoTsf54GAwoP
0g6145Id7Jvsw0WIfo+PJ2eQNXAfh624I9dNs2ukRUPhpEY27m37eJo3ibTOX0/KSA8PAlhjOKRe
HQwWRj7G5h1drHjAh4qL55RLKclWkB5wCPIcb5YJVsNPrZ2M0EYzWOf+erV+FgevSMvu5RfcQkah
WecIAPHGuYjSj39P98YEAMPsLXIvWfuBhOLT1sinPSDUsmstlcMO5ggPw1ClBCZyA+vbEifIewqv
C+pVv+mpXrto9Ggb9wEe6x+SnHY/Bkytn16cshdQ6lZzrArpD1TFKrbbzZTMHMul++5DWmCh9WV5
r3TNcgVdHkf8lQ1kGKSs0Epwln33W8XVqas+ctVyOGCAOeLoaUndD1NSdgKlVnN85SHsn/fKxw7/
k1GHHckRqiLX26FwxGInd8aJOainEpSslA8tri2AwYZ4aCWtHW4z0bRNJv2XxTWy5dxfrYPtl4Lr
KDL19VoGeZgl3Vl3QqCHZHgrwEZcWRdfgCyw67alGhS2ucYLTF/z7HqAWcbixmL4+9I/llXxZLVC
ics/qvgI8UBPhZbVdKcZIF7DE/vTlaoJ0WW/QAk3y/qx77rZBmJC4PSg/TK4BNncsDvJfDxgaSTC
mmdXcVQLn4k97VeYhHPy68o0xs9vsjX33RQVD4kDFMP5OnSl3CFS51orTiBiAOBqV0DfoB6jP1Rf
tIlUCeDy4uBZRG09QcJHq4HPuQHfeFx4sBBkuIG6EqsP11Qn7buEulSJ3ZYVaRHrSLBGQYxG/NEd
ceEPCfPAhASlpoOrrz0fViB+hp2aCOwutvpb4KPg/5e5LfRySYneNomvdYEYN5By6PKxuqwftWop
Y7NTq3A5EPLOYKt4hnKp25lAz9HYcSk048N+Y8LN6xNr7XqJxkbOaeFnkw5JjfVPkJQWanmaBHP1
jbfl0rNNnhFEAlGhDaH7gP5zA9o1Xc9HMlSnOoltVfxgUrlHmgTJVpeGDd+3KU2gnVJQcCGX8hBA
bfJw3FMgsjPYkbf5lSsiF8jBN40Zha3uOOy6hzpNgL5wYYzuHTdwusAuM45QDN2SdE/Nat2gYMKx
Si6ICocxFgg/RRqJMKErLjCr9Ay8S6Wl6XonI03nZQJYCWCKGWsF9Z6HGg7a8CkotAonGDr3G5Te
uJlO1cusRAjVyAKlZ4cu8V+n6X0fw0RP8Ze9TO/APt/UU7WOh1Y6PQlOggw7eo8FddIQ6zgm6SGd
EMoSsbdUmbl4zI8CC6JvSJ3GwqjmoEmQi0p1zhEwKRJS8FMLm0EkxqLNQwn/4u/aqntGW/qT5hif
YuvEAVZAbjv1nOXitq5t+NBsVKbh2nmGSpfamHgE9YOtDyysywiobQEEjwwD8M/sQUaTQh0MKRCe
oOPWfoZj2NrZ2JN6LN9gdNd2cr902eMX+SIe0RfK99IkfRki12vuKqwvpQE5qLu3Z5y4zKQlGTkJ
CL0q72cjA9DeHFFDu2UIsNJ3Osz3jPw9EIZ91MheXx4Q7lc4XD5+lFtEtGncuXcW9oXIY149po64
tzNYrKXO8O8YY3Y963wlvDWrWNch/uXlOle84ooJGs4xq7ks+O3Nw0/fn4JWo3ZanXjcvB4mqkow
kcIk0a3h4gINoiQqY8M2AM719TZGZHo/842yWz7JMPnaUXoCmHUgD8lYoP/K5MNahzG+77U59bEd
MLrssxDfBlqKeTtCkquz7BxswuNbjpAA7LvlATcMVKeTBMejECsvbYzpZxL5zqUZGCJLnnLpBwgP
n6loDINaZcF284+hVLlMB29HRUAIeoJWMv8G4oKq3Lp2BX+U7PqEy2Eyz/YMz7OAqaIIbFLbFSnw
Wmrg+IzFX2lhoM76usmYyGclhM5FEb0ltJqiF+y546xofbdJYPC4OWCAnjH8TiB9K83dT7kNE+hn
ARNOJiylUQLWkQSxuk3S+T4+pEgO8kWl9reiOQ4OVQZOyYoapK44e0R+vzEWU/jgDNUyIbFHmeCh
lmrjsWOzbD8ib8WQcxOMyAPPinfPlDAVZ6KoRaP9qVGjuLUll9MexX2HyDiHzx2bIqqLP1XkulKP
/MJndRJ4zUqdOgf9iBL8xS6X6m7+p08bRJzr3mbKJ1jbIztacAXjmKJLOU6QGQaB+cKOMBkocyk8
ozdXGo2hlW0KwJzON3YJk/oVZX6BbBOqfGYovD3msLa2bzGIfI1bul2Ayxss1Xr1tAH+ofy0TuvK
LuiaT93FnAVkmFOoE0LnSBQii2g1lrYyBikGTrdVXEh42Jkw9Xs7XzOBNS3OlbNpdEVdPxeX6o/o
w5f5ThU7zJbRBZFz4sG2GwvlyLpPY0SeYKSFnUsNRtHpzzUG0cjsfDqxDQgYiiiwO9XMcwTDHGrJ
854hYsHcfL+X5/xG+8KUk/dyYWqVXTzWkGhPHchBJGnt9S+AZHSq/cv0/uynhb0GGx4fq6QEJ5yk
IjbeARnC9phB0zDKfyFk7Er92oMRhpRr5jFXZxIrjvQcEH1RPrzHSFYR/KAY6oewoWKPCuABp6pV
+9+Kyk0glyqc7gEWj8q9nMKSL9JXTXMoRlFSoMR06Rx9W7PuGI69ITFHssGyQJr5ognpd3NyEcKx
MR+07k14IBi1VtO7wzgIDSanQchFdNY2+oNZ6AZpX05O54bM1Dr5qEIdwXDtmnr8impCTNce83V5
pYonQXUHFOZUBiod6b8v1I5j6y4vOAGtbGERad+qQ2P6akT7cygNHSVlne2+6V1jvttjeEoCRcgn
aXAW9Us9+mjp9esfSx/2rRHM8iE5cdp0zFAOnTd9wHlZ2kwHrERfKT2ubf3Epkm/R5JARpoiXnuZ
ALtQoxnJdrwd08qSQ5xQe5xsIWsO+AMGYxq7P9r8JlXNfGuH+T6UxnpYqcJwiXVNZtVIe4JLvY1d
79gSY9NSFWpfTBEObwlvNSXanMwX28/Uovav3Ff1fF4VLy9g31yFKd20b89Jh88FFdFrIUaWoOSi
0qJumyi/TOyhON0N4Pn0RXpCxFXEzxBdWTfmt0BVEBSrPZVGdkYzU95R+6dufs/eHCtqTr8b7wz6
W0cVSAAYR06pHnOQSaNPWTjBFJDtc1K+lCC1hX9eW7O1/xBEtxbOradH3FqPWZaGWAoS4a6vF8iQ
ak6VKnUVNFdUaIfzUHGdNEiOi9El7w/A27jsBjvGFnbp13a4LS4DgR3Ygdz68Qp5bDKNPlDlEHLv
uvwEOKFGVlLIyur0AqHXs0LWLrXrB+0akpycFk7jxu7t8KJxpFkAK15WeowCRAlh/Me1F0TUNBg+
0KjV5DsdR+hAMb0NmGssdPhE3yki8ULJIDXsgum2xICS+MsoJIaRNi+dicfps2pc4PvyT3uELlwK
bi+yPPbriqS/gZSxjgmeO/RR7ESnasXeUBUts5ndi24rcnZyJt1aE6uFTAomK3sAw5lRVq/Lsw/D
p2weCsAGgHsp5M51E2/N64PME7Lo8y8fx4HP2KVc6p+ZBv+Ut6W6mtkfcu1/v4jWCMrNVHGB7JUZ
yXBAH2QZ5KiW4qgq9ClOrPeZIrG1OPxQ+3smrpRXo+BWDUdacnWGBtJYF+qpXXRctkjPV1hnYLM/
guXa++6UvAoukKr8s3Jmkehcpd57kRP3Hl+5NfDtHCA7YsJUlaU42rCys8uLIxsv75Q/4HNIVFJB
xg5k7qA8qXA8YzSVdtH86HCc5/bZMBSRie75Iie4D+7/VAGqe8CbCRf+IAoJxR3ZGARbAaNzDlUZ
aAJPoA5UoiC+dJr4MAG+u61LdztWT1AGPDeWctibNlMyrG4CFoglra1Magyqyh0GgRHiRZjlapWj
WqgeWQGQt8PMvdvEtOL7hW5cBQGqbhRTSczcyDkhptYBAK6BfoSCU3mx/zg4niGhdLN4o09ZzclJ
tdwkmhM0KDZV/6I0VoqtvZODDc9zQkCMZoFEbG1gKkl/gRCLDbupEDYC8XLYpm/uHvJzFoWqw1dO
klZydDrq9OZ6an1AtOTuFMfLYxnIyXK/qhKCC5ARgwLaQvGq3E3cUm/Dm6o/JHznZhy1V9FD5z2e
ABpBL6kTCjMm6P9cWWee70hn3bYCo7srhDsEp7NAlqh6s3SDHoDIMBFITOjqqRRCsLNeecspvzIE
j8IxEqkJwdooeRULMEiWOkLKHP4V05aPDngP+k86QCRJ8gzD9I/7It6bR9QuabI8SiY6Art3ev8Y
4RcOdS1kUbDAQb/NEKDsMaDyW9nRhk+ONuU+urqt5s4g4YDcCpOP2DIm0uOFWMyq0+Q8OXi3fxT+
qYzzB91sGX/jv4MCASrbUJMlIfTC8On83ggkXpZwCQYvFumPPb7hWXeD5wuWwAiS+gRhnfB6GFcZ
Gliip3LgFszoBGiOGey9xUro6RHe8cPaM1Q+jPHEzO7y5pJltwRzBKc4wiAjAv0DkynLSFiiiDKK
FcsGiej73ORcYXzToQKV2DohesVuuNmQGQlkToLxkzuO0CeMoc9bcYi2rJxL4N+Vhy0vJomOpwiz
pb7CcSw0Q2H7op9XoD0+UhnzVikD1Mhq/O7A2xOHd/tAgC/qDQrKp+ykZGAH0dhiEgI1Ja5s4R5G
9zgY5sYkWqBWxjMe/nK0PL/Iaa54ofJxeWjjUiOf70LH/OCHYB8hm/ggy9kT9CFB7p8uX3BhXQAz
yrfj7KFStWS0pElwigWbMqaNlBhW+wLZPIxdHXY00dfWmT7k4c6v6VEat/6Zc+TzA08jkFsXgdxT
wsL3J0cTS3pYJwe8UzcOpwRDurYJ4UPmDKyBeoKgFpq308zTKp3i1+d4a81EJCQ7OCcZ6cWQ+yv/
Uw/ovFT6h9zS0rVqzP0IgWln53YMwLjlFIV5T8P+mwXEPxH9rELSRWks0Ywj66EMsCSc2txghsqI
eOwk0T0LxCz+d7pnBmpEfZ/RTZer+BQucmt2nUNKhg+sjnpctd0X1WeuLyG6JxTWlZJU5fztVfas
koDe45KjfnKvfrIS+z+1aekHUqfTDM5l8+yr22oFynxKVuubpKPgj7ZlLdFpP7okXL6u88eiJaus
YZk5mVC2Am2ifXcWD9dngA0Qg0w0xRuaylW0BNjvSlIy6LH7im8hBFRlSHjuFtx3R/3zvWS+p+YV
ohAtRmX2vzqEW8LeS248IeecY9SaaQv9K6Vewd0mP56Mx8JnA+ngaVZ2wVG9V0OchBw8m92U8gHr
ImasMyMW6yf8nJpawxc3tLiY2Lm7i8O9zLfsudv98JsHxmsahFZZ+AfCUu5FvZh44AopAfT4KKdV
Apv00fLN7mC2avwG/X8aMfmYPmrsDIwIoA30sYDJvaHUWRYj6qk+W5OYTDUQqSwO4frtAu3PeYrG
KjXYnIMvg6nhBX6jXy3wSIR69zUhF764eQsaR2+06dJzVSyxgpS+R4UmxNJR03gNenm1WG20o2FN
oVFMfXAHvr2HHyGpewQ20lLJ2371SzFfwLJPeiL6Ga1uG/3IHrWNS+mO8c0CamYzuv/NwwH2QKFs
jR9Wv05ogxR4rydyhFnznMMIUg+8D462FxiDbJN7feE9gidfrxmz2B707L1KiA/q/Cp7kl+G0D+r
qdt7T4ES6DknvBJFw+7RiDLrcL5goYDqJSr/wR/DEni9tR8vlO7DAMh+ImanUyREwu5Lci+FUZPc
U+RtDHYEtkGzcUQV+2e4B4/DaBsHqGH+JKopxR9waCF2syoyBVMQWrj5j31E2KKF9yNSIwwtrOAa
dIalcfhMYE5VGyRnyTvi1zxNngV6FzuoNeMaVb2FRtASbSQJwUKz5TtT2ans3PCpUd4bKP3o9vjx
RZBRpiaKhQaQvHSTkyr3cMKG+B9B5ocwRJinPryouhy1O3hWxMffuKOiU1IpwTKfTKf2xX15UiPc
tVk5Tk9IwBG5ZwV+wsjSfs1BNaP2DXui1/HGJCZw/a/6SMiCcZuZ3R7Juu9OHamZggG4xzW6OFLy
XQ8uA4sF2AelkVmsq4CJgDF4O1WYlD1xT48WIjpa6XhuMgw6Au1wkGqC/KWExmJc1GI2VF8r7Pna
5Qq4xcHrGb49tIsNodFfTF7PSnBWjz150Hky86E9HJTak0UOBCo7EAENilieK++SgLhYPm7R8FjK
9VecFUSz9udabqMrLDGRJTM8LyTvrCxpTxf5qKjoivbmoCLki0o545JW/eZoJexwkFM0nJb5cqR0
2dKf1js+53NNIi6+4CiB7yuvFHUiJJfbXZ610TMTILiIaDANqZxWBduDWUAcUOxfMBYvU2Mn6VTH
5SF6SFMogmp7jVnX+qnRsCMLpDjEElqps1/WrUB1bjv9LRUFpvTl2xJ9AAjYuYxYm+fXo9o1cTy4
h6z6jS5quylKfp6C+y7ItstqVFUKaBz1stHWV2oo3maOQUP530aBJWmxuiRvJLO5C+Z4mpZa9uFi
2exT7Suu7PUTsyWYHSf/1iuwFA24pyPW4zWQ1j3vjRDK6TMOMdjlFavM4uPwW4l/vdCdrBOQNh9K
kAoCJCAG421m7a3HuKvAATOOaLTsmF7R/OnbTdsUYtmrCRqXqWTrIJRIJf0epShd/PhPsrmU+kBg
lHSSMqAuxYx86MraXCqpU4j3Np8uZJUO3fE8TDlZ0YYJPa4EdtGbh7DLm8+CovdGV6ryHOIW2Ewr
KujoOe/jgFY4/eNoMGpVBv3a2lyw2e9hbzI4HAHhSyGdzOm3IU10yrs3zp8yFnljI+/xNKerPQ9e
92J1AE1SfW9aiSx5sfgVPtdXSHHh0W0oCUDwmXg6w0HPsjXjSPB98jbFn1OnBK/VNbH7JXqIR+tO
dBsZEk42qTXepA5/D0FiRx7hmxzbjv9C5F2i4oCZTsLLTy3GLM86kWKfnkDd8KFkkK97AkBgBTfH
YrKyQynZzZqXFJuodOuck8jZNOd6bF+gnCa9gygyJTO11UZ2lNyf4HWL8xKok7AhOdxIdldzAh/S
rpg3v2DkDtX2xJFgETMFQcawB31UW8zfejnhim3LPGnRvF4TdqUWA6Dm/gVPXVKriR2DegkjPhi4
5nIs+7emgwd9aVnx8nVHKi8GPeUpJMY+owaodvZ+IVs4czNsjL4oW+dDf4MqNmZLlLbhVxqXoH8x
sN87LzrElR7x5FB0/6s4uJutZAZU7FQOLplUl5c8j9Zhedw8pGJrCUjMBBaoDousY5Des6PWtZTh
sO2iq3g0Ptib9adUDi8FhEeRwlKCxgZQ/FFtsTIVc6E0PFscyM5SpW8uQ9LSe+4PDdSyoNl1LIUs
MeDxcE6SUL7680xAIpqx1BmiEU6Zpmu/qsIRoWV/igITZfwDcVcjugaYQwkzrSb6icV1UBgsZYfu
P+0T4T2bDOBLbCnkNe7Surp0kjf+QY58OOI1B0tWa72NKVrax7iNe/wEekLkWlr2QDARJFAx20p3
Ft2by6bQqDVIUiydTgm2DOWQNbAGmjYSjXA+jxAAj8Bt+R+Dpi0/VSgmBtpeDZ7VvlC8qb3IBROe
uEsP8WXvxDizCBnUHAfIpaibZeCeeHt91kaSmsSmhphg1ead2JwbxTjj69oO3rhcmmgigHNkrOHu
ZAqrgwgyiIl6FFceABNqeRm4nGqzIqD2BtRzYXboIhyDonXTrm3x4TOp/4riGpbH/NSHd+Y3dS5C
k44EInNLV7hnweAi4B3gjeEX1prV80J9b5UhSfmn8HcQvZnheqqwBRJUJzuzRI8dpHaWT2/vkoJ9
7FejqYuQe7c6ddBrKATmQ6glB5HG2dO1GfKoCRImup8wyeCWcCVC7lLWj9KvBrhwBCisSlvvJD5l
5be6sxFna2BzFok7c78vlQRrRWFHq+CQGdLd1gs3DkzJ6rR9T5KzZZdjSKJLhn0ZC9cHzmdGMkhh
ZxlMlXG73bWeUTSVIij7pyYVbhqkLO4bcurW9Kef5STHDOgCCr9n9b0WXd9jvidtxf+veKp46j2B
P1Wf8J9iAtNSLapABDu2xO0COkc6zaGADbBxfrmlqG1Gmg3yFNlmjUzJKOR580LDu5xaBdWLPsuV
oZv2vk6zYQnO3oTzpepoISbt2VACSSBpdvh5bX+r1crMP4XB8tygC00eZWrwA+1zvouhuR+JzSWU
AcpHRYuGAvylSL/T5wwaNfDw46N5JAialsEYZvz4eVtiaTki61owEkOBX7hkvZ7HX6iUBRhKa0n5
1mjqxRPrA//q+7w1pJnWajLe62OhoZaX1b8XdIY8LfLyH1sWLYXlDxmXGIjdHsTdBrisfPzeggso
KkT5BFqucTK9QNfhmxDCjydgFzyRx2Ry3ljL3BfE22l05hu0NWegrFr8p+yR/CAPhK2JLjsuaNtf
jtoVKma+9Nz4F9U/J4WWcrGFiRI8UxXe7LOrbfWMFU+lXtPB+Nur0pR4YNnoCIgTs7too21TtGQp
NtGxBxsPXShNDuLiOA9iz+vVpP5NZa3GQXIAU/hwMMzj2GMLuMs9ywXeGgIr2LZnyMPahd/vWJXv
hBwgL+KVvEAf/EJsHxCnw9p0P7eDBuJ0G4r3rMKFMayERWnsGRe91o/y0SIGfS07v4XBBwgHbdLP
KQHY14vHTfljYSJagT/6pjuCiRxZmViiZlNmpx8lilFZ+KiFJdIZNSkV2g0rJMTIblz4/ArYY9Gx
RF2IIy4SxEOxBG9VgphysYbmq3dXq5JxoXCIfxdriS5k8kSf2r/6tUFwGjD26iQANgGLOs6yX0Kr
qbdgRNaKU4xx1S1PyHFpevIBDJQ6pFqbkDxoWvnCAdlkmqrzbQGJM+RfLTLxWFos6RC/N8uVInlt
hxsZmPHABr4GXygXS1lg6o3LiqTAqUJmi4Ea15oJE9iw/snrPCbujJvD22/Gtb9CUjSmBy3Mi1dF
OBlMrWUKmeQUo8/0dv/dKKDszhOhbkWyYvc8kkfpkAoziAaeDWguOqdGlpFv2sxLYGpZVdvOoGJN
19QYkQ+WI/b/kgP0FG68fTLGUFqgT/udFVnY/X+L4SJJsVnPICw2BdKSo1rhet3gjp1ZIi6MKX7/
y6RO8jHMLRuh66cY6+A+06V5RnD1YvliXJqN4DYVBMRCWSV+3RCKggLaHIRhmT2erkFw1h0s65ee
tCxv7xKgADxBhr15I1urzOTuQQl3bdhqgcuDw8A+1utkBlUhQqq8PObgxMb11Fdie5d6eMhzYncN
LFKUy+vhjtupRT1OIweJl6Gwof6HYEraAMyHGVhZ+UkkjP0u6pgDDBwJKcRCYlnF9xFNnTPt6Ne4
sGoUyz3xznN053GwMwi7FmKCBX/5vGnHJ83qeLzZMMUmhQG8uEUpZbjohlmoapFYQcD9xoAcDC5t
Tuu33Gt1Zv5Qbp5vwZc93pjhmJlxGUN6/fbsSuXo4ObQgjfy56XIyeiwPx+kcaC6KFansnEhLbUo
j0ydoT4i/LCeleDLFccXBCvAcJoAjn0M43J1R0rjJjmsl/+DoSNWUDQL0TrsZcmY6lfIj1VqOvnB
5q+KhnNBjmqjokVU1nSxb6cJcLBmxRxIlybIRiWUMdsxCNQ/B0MV6ieK0OVG8uO0RSigdvEcfmI9
T4VvQc42PWHYEqqtQlAqJsgXYaOOJe32X8502659l+0x7FPiO+994AK6+pf41cVUQyOjAmkLg8yY
hr13tJoFd14UYtaZbMho91h0CIeBx05MygIf1M6r1/wtn4LeW8tGYizb3Pa/je7Y31/RWNzWav9v
krYZ/VBEPuVHB7cV7PlLVlXNBeSqeMqm9IrzeAxRp0s82y3ThfNn8bmh2nzXWRGvGnBpapx/z66z
9zBeJMjsdzGFZKbHaR+kh7XO/U6Zc+MSEOSjgSCZYoxpxiu3exwOGucBRBW55I+VWuMfWAeXU3o+
frFrNK48KQlZeCsMAiR8VlAQaDe5Pub8xDE1BZZbe1dCGkkMJMSgHgNzzGClnf3C8Emq40EZlIQK
XLGDaE1T0CPsIxfLRQecx7KnVrsqcXNeI+utIPedEmRGboHVqmlCKqnKgzKznZCacfkzI02aRLmz
UtW7xqo9bqBZbwss08aZo/DUm4pzTyjL0I5NQ/jCd7HcIlCUmx07a5JLly1oKgeaqnj/PEhsEqSM
tXys2OryU+cXwcdnPM0/3ii0ylc+uyXDsjaoemBvaIgHzEqmbaOk17Rc1Xkc93S9nByW8uonrzvJ
wDx0gG6e+2Znb5P9w/t9rx00CPUCk0FmZefzqGSznD6pV22Zk+Ol0Vn48DRoMsVdhZvS0YuFyUGd
quEE+jxV3eUzkhcoVKU/URho/d5+CihCinN35mko184AFjyKZ+3Kt5fkkdG9BVZwQ0Tu6yZebzlY
qDbxPEoTne26qzKFQN7KIjoO0bWiN6fAkKYpbYS59mYjSglIAfhAmtxTOSlhbXS8Bq2VtK8ktCR1
wfXRHGVURcmZn/5YDSUVsGp9gWPQV7jg2qj7Gc4qcO3PVpV5UXl+5at49l61YFojcarVbeYxtWqM
gJjJrOYUk0LrDEqduVROLFZOuWhLOtdA2j1iR4tXfHfRylbRd3HTAzI7PzKREzYaugLCE2ncuJhW
FFmvI82ydT/tuh5PASR8ry5MEmzAQxyq6ogHgQ60VPTyP0sGI4ns+dUhvU5HKP/AF4atqtmNZyJL
UVTAljkRZVm3ZhoJGSajJchak1zjDBf4rrY+Y0ayg9YsPxPVkMrhQc0VWr0HQfogrlqqGB1wGlcw
prEvhghX4R3K0NgUqO/rhJrqXcIAFD8D5L7VvczeZbBFiTiSzebbfdMsGy+FrqXrJeMt6/Zgs9RO
iZu2pX1yfgWcJd3QopsIWnBe7Voircf1BN4R+E8lcoJMA4SKpoIMGwbhJcr6LsgeyKAwqEMn3Bzr
czKhJTAsEQnnJWdZh71PiUmLWr6f9ungREhdjTlUKhnOZdNwFFzRBNpSu3Vjwg37peuplJNesYLk
lSyji6e3VKnAv7uPCql1ccHTqnBoDbF1SoTj1QDtMU5n5I7gYuLtPZ4ChE5uLkLP4+Jv83d8X9h4
oKRE04ZYbnTzly3L9PRjQ+M6f5oTgDQ83u2h7FGkn9YOLE3rWBdqIwIYTbh04MFZIUSPwMMAVS8n
pR6pDJjHGyJjSSnDIulWxH1nWwWcIFyERjntAXv1NQKlADFeqNVYAJJH7qQ1+xfynzvVAE0tlKbT
4ovOoZhUiXeEr+oD8mwqC+1Hq8XBGAUtJzal3o5MgF/QRPHSkRh1xfXpcRxXZKDovjVPsPtbkRTw
NaTtmOKiCFLobDj6NiBUzR6yOsG1sgwO0ItmGj7tO0gsOTIHv/uebGvSIceCw2NKuZyKxWl7RCyw
WI410oATGQYWyNipJJ9Bpokdzf1yAlUBukd7te12CUnETyHrbKBABKbvw+vu0EKE75T1NiwV3rfM
LYDTmvvvcj0yZE7lopst5iUPbj4u6gPSQNNOsu851torRllK7EX8nfEgLlFrt1fvk5MUBrl9an3B
eTmg7+Br39/Fn11eor4+4efwlwrMjDzezcn2I9ecfojeeqgZmY/mKSIQCgBEUfrGjWBtQTX32scB
qprcd3Oi+mD2acDtvRaVA+Vt6nCX/sF6QGmT2I4VT2anEgaHzBNu8Gf08JjjDv/ph9D7lvOpBVIy
0iq9JEyA/meWfNW9iQ6ow/1uUtCm5JBCNqrIYhtwDlFL4Y/SAp0a0ew4PfLWIDJyRhTUuZnBggeM
to3JoyBRQkT7gfQaHs8tqCP0G/KijRFVn1MOXiNb99KeaGBnQy27J6ZTLel7catozj5xwbzubtNF
XNPHAEmgXwZZP73E2VUsF8Vv+WI+F+7+VTRiAY3ERYqkfGb31GVLp1jXHNyJSvrlBcgz4t9tXi10
x5XoYsegbiSnUWN5DPkXJmfEakprAqH1A6dmC6CALIV/glge9PhIW4zJS4m48T02eThDLmZ8E5no
wKSH/nf0t2R1M0WKlpi0J85lHXThPfkbsUjOHRqi+S0kkofLCdo6DHy5QKw28CSch4mMDKxie6N6
HzEbq9mpNlZ8iLRTxWDoj1xXv38P2VMslc3IiEJr5Rfodu02jKh6DbQos+N4S+ZQSRMbfoR7f21Y
PsY7INJn82bV2AGP5VpvTd1KbQr5geZeDJ7D9wYnpOT3FYKPNFFyXOtdyC/h2UlRP4iIRPnKmLkz
t3sN2i60E/h3Db7V6ZP1eLsirROv8sbpXKxKBGLo4vQLRXB73+aThVz6SLjCck03uKELthrAVlAA
pyo+qBVlqknret+ZdXeVAA8wQavbEya6DnVX87s1WBd3OvPUWOmkndTyDwIz0yACbtWcPy1Ce3Fc
ggLw7AYNo+wZFKZtMiPljanaFDkDL9iGo6Oc/EajJbzGGFScEU8pE9ag22808LLpu8rd47kR4317
MRhZExXL97+tg5XXtGVymdL/AjuphdLC49CB/u9AvLqbujmb0ndzKRNUGg+yUz7W5ayFTL+TPnTN
YsbpZuJGScqiLJLpNfRsPK4Od3JJzHRhaw8tRD/c5E+43cmNAvDj/quG6JOd2u69Ez9wUs/h1ocU
AJOhQoThvqw/rxNgjoJqEk0MaNSySNpV+iqo+YFU7ZoYO5D9dTmi40szT1CouLwY/2y1N5mWM6qE
17hLn0CRNCQotCcI9gFJ564awKRUgApRBWHdma15gkPk/j/hB0ixx3mqSVpIISvc8xJs9ocxRz3m
qXaYgRJz8ubkZ4C05otZjKJfYAXAnt9EpuxoK6kyUXhxxWjAsdeHNbaJXmbdWuYBPvSjBZdU6AEh
cHUFiKblL3KkXS8fe0ml6l+3jZ8hDb+xGG3mr2kLeKbH8DdRqzxYMVzG/mi+Vn4QGaa+skfsDoTF
a3A6G40Z40wd6eSAguVs/CrPrvrirZIWS5TZvM0wWfYJ5rsA5NZqBsQ0p4pRi7FGXKIQFXok9Uyw
o3zboo/N30EVw1i+IPlRk75OA2RjWhSHY8zr7AEXhd7Ug6EhrqZxBLWzudBEQBigYhnwtyxw7HlS
Xmb0BG33LvHeSpUjLkWr3bEvt/TnCxn4qMoPpul0XR6a9a0t31K8i6BLhJ1/d1SOW3XSVpZ8abnN
9oR82LT/vSoRkgLfbyIJIYNKkHeDJYnkAWnB03Wo6c5N6PNiFnxMpcBPH1f1FCOfdAAY7xtCRoJu
cUofFtAqAl+nBZXNF6bnJZTFX6qPxPgMHrcNweiescmwlYXgmx2k9yGYJ1voOjsZwegjB3krv75y
9Miwo/mw6E2qKg0Z/BvsHEkK23JYV3it+z4k2CTzaJKhcYCU485DOkGfrLHKHHuRoCOL2HD4QOlR
nLX0mCRZ+nIXFswn4GCv3toiqDEKRaKWo1mCivyXdJ/kOcTlUdic+MiCv1+FkU4gxAbnKtxia2o5
jbP62RFAnkC7nVxw1HaqA8z7wYNXobbnJE9AFTjkos8pkODvzd3/cSJSapg+sOjZ/U7oF4CBk732
7xZ6KItHBAITwfmwkpv/DkdYuAGVTdnAwoYEoydpT82n/dd5szWsLYoHhpXUSLQ+c48Cu76fSivM
Bpyoh5WjmoTygwtNHt50G4c3YTf4PiVoq+OiKTS21qa11vetvolGLmkrGVRflfcIO8JF4hVu8KB6
BtZ85o38RDm+6o26IYfhwh1A255dKhii/1fSEbDZweLsAnfx/0JOknC94p/IxmaoE6cbsUf3HoMm
UVlYPDNVBa92ehBS7Df4VHegZJqBb52B90HrqjJ+zMuC/8o/fYgIXP1+E22XrvDVXqin8Z8wsU4y
Pisu9FDLv7umZhOTy5RRwG/7by6foAQ5Q6hECOgtY349CdbJkKzeLtihS7/coSUayhYQvKnaxPYC
xcntur1u5g7FprxxZlDAcykucyS9vDnnJ+kAlB6HWiDleRhV/EYtorTAlKCzb1KZCNWwTM+SbQcI
7F+9LTaf0q3KIVT7A6+QV9teguSIhmNbXrdh1NB30r4BmSAeoT4sARFCWJwqpgQhVc5pxgAqjAVv
K6mLrhwN4rhzZFjRrWiOukVnu19tNJH/QreswHk1mgpFsaEVri5o76dK+q81JLgGw2el0gJMm2iQ
cN1HB9SiAYVfJf2/nGpij33zlvh5sMcoUHoqqzNzAFRzs65rCduDK4BEV317T5duCT+6JOaHB18/
qX9P7LC6Z9TEzO+I9tejqu2LqOdXOkrqW0vAGvsXGlR8b8Q/prAR7sC8NSmco8QRgCEnuc2P4sgW
N+65P0DEiS/RcqNwUWSrJlIhjgG3PjS2ODonVPLU5WUIODnddoslsI3ix+NQ9QEQ0S+PGc2M5/nb
CeNTsuykXqE5B1tiW3cEufkYNI68rGFwCV3AkAaWLiC5TbSl2vVgqiw9Nmj6J3V4PkdyRf+XgtK1
m/ztdBWeTWco4pjz7MPkq1SE903OHwynf1+0P7F3AdgHRo49D88L+AnUDplKUkEUrXVPf1LBMru7
+eJ1ECDPeF3VvwrNrIViVNOTt4H3JR6sdhn4A7EQUge3A2fAdXfbodnVRTA7/UEnEbFOM81L6Ukz
OV4tSGNPbpWWjyDT1PaIOWTAqSszNKW7LgLwCcM/U6JElvSzcYVsC2Y3FKVQ1qbwLmvJih/bIwXD
OC53POseSOknUAVC0lxTcMi0B4z3Ts/e60ZJT4mLxF6gUc2nbr63brKBYS56n1VuJzhPRBaOFLg=
`protect end_protected
