`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Y65/MFXWhhADwOVv/M4+o8eaVO22scaJrgCxDXOByJVk85241NyhfA5m0IyE4wQJmggZhYij4hhT
+3kX1z/WLw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZkenUivUwQ4WI4NH09hs8kGW6MMq4uVGfw/NDOOC+R14rbma7ZeAsZ3KqSxlJgje8I/XUuGZog+Q
BqQgUXa+ZgnYgmCAp0+g5H/YK8jcG2T9DuF4eM1S2TWLZfAaJ6+Oih5mPKEgnSN33pe2nuPG/tCZ
WXp1OZFZ+RB/28BEUq0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KfYMeFs5V78k6nww/KOz0zj+63zNb4UOtAYickTFxZ+X2Bnwv4bsMA1cXnQyk4SRjC7e1wBUUIR4
UfTpnVYzTQ8JpcBUueX6sU4fNn+O7u+hXQUfZAI3YMihyTW0Qh5TEK+Y0Uey1NL7nPsKoI1AWQ70
umGRh89sWKiT/oKyLtcRew/ZbNUPpJUMKp9lrijWopqWCeA5ZLFHUV2A31jPWLd6eOES4Ksq6rju
hbFRC+a1t8uoCoTa2PZzl+q595bGHK6L3br1Ee+Q4vWmyblGzhWm0BAImBBFo7rXmogRR9sSFa7r
Pn0ukX6kc6eftG4ZTJ+XUDMCau0/outNM4zjsw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a1bFcIkZo4zPJvMJud4vhE1uFKNbhylkuzUR4O2EkGwLrE17fGyp+MqRG7r5NXGWXZuU9WK/9Gjk
0rdtGmDcrDBvQvdIzWLM9suFKzfFzhT8kOH8hlb3G83f3ynzmwpzUUgKGmf7tSHA7vQcdXCyq3MY
kFp+tB7AzWsmU5Ifzj0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wS7l1EcN9oGmeOh2wHa8aGY4hTUVFraqFIuVxqm0oqEK6gJ2RQD6ljT4vhdDVHw5uWV27xjMC6Nq
3j6hLI5z6lDKEjZm6dNt32pWA6dw7FadASbVwuaCyLQwHr+jXMBETZB6CFmopdxOWk0tjAmuNT8S
6rrK+f1fNYptaPKfOjH2eU7LJItbPRRhiA0sHPOwWzftgFEnTC3GPMw/GNmRFIVoNJWdXxbY2F5X
9jIl0f1Yz91j0MvUjp93SfLG+NrxinVmKZNyCPJxurpHvwOuxUesjDXLOc7aaF+A/2LfTEk2hzWV
MhiTwFpPJdDm6LIJJhpCOu3SBVA2U3JHuMoe/w==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BfNd2bDGBtVeSwbNHF20kdZMav8Ejx5EwGOiOgAGrQhSyAHpuGt/EXA501iAxaGv2XOVUgjVCInS
6ZqAXdnq8jYBca6BFfB75y3N2lAKe2aXiu1WWsOyb6BrcIyOQojTYsLNE9LwQktidMkkFBM7XJIj
HYLWwK7vKg9moWzSIe96UK+ymfjAGVJFjMRtSVMdHAbKrQWC/dZH4cYbRVC4BDkNzqV37knm0PDx
L+DaSzp61qE/otP3FteBgrxdQ1xkZWWq18DuN4gKD+tcxw79LCeiimII2/2/qAe3L7sYLPUZMih1
XflOAcTbAMQkdolvxpm7dxjneu28qIJPdA8CKQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 637968)
`protect data_block
ZB9h2BkRgORVefM+y5dAkYxHKEEqSyrkVFeVxrdKMekH/2H5Y+c1HxJ53TxI6Z09wFD8JGDD9DwT
3fsecDj/8c5aNyYSyU7mg46rEunkyCtuYK8KHV3A2pzVGUHXjpoVXp0kc/kTgG9/MfWopGPDSWsV
o4s/v7CM0U0az+vxPDdzCwpazYIq5QvZ3I1kWFuALgK9d5ssH0X4bY+/q7v2cB7pbiI+50fcWM+z
mZ97sq5E4Opnzg8Tm2DY+PvYoJ46pU+rEChaSKybUL1/0H/zZlWNs1rEECMTQNgpLD1F4OrlOWe2
AkIZve/gzt7S8fPayMSfMfDkn/IyeKbxqi6TXkhYlYO38rNh3p5wGXaiTWCFWmoTQWEe1xKh+alo
VHYCIxWfGjZ6rm8B8daxBj5R+KDpe+5i9O4wPsTMOB1lhVV+gRxbG5gQXdT1wTWGwx9shERmSj49
hdj4taDTD/g1tuAbY7U5xTZ1qk3XSlZLjYE+AvAYpT3nwo0Fzq8DDcdqaB4idnbpnemvlA3xORCx
xyHHV9Qs177PUrlhP95nbHhpya4wMyLFu/4mjxLhe+AIY8Cpo16nst5TyQetkdFqr/CxzjnTXGdf
pXgjvexVq7lAcSdDt4j2C1lFDPy+WuKjwWezjYqaI+7awsIjR4Nju7iRqhyPWol3km83FKjQQNrQ
860KKwtq4eFNohd/9Uy4apqjol7F0EViyhUICsQ6dQ5Uaf1eMwGn+LwtfquvIgCp6tPB83r+fiBd
Lkctl/S0y9SDD+zKcxEM9KXH+Ei+/kl9L5hr70flns041RwezZY7dgx9VRSVGkQZ/uv5CgSy53go
StU9VVdZSpXmXEdXl/CNw21OIKWENhhcI/TfoxVfC2tCrmbvSMALNha4mRNZ6C0NhuHhVDkmCuh6
kiJVfMAr7oniWau6SZYua7pIGtThz9j8zvuLkDG3B2UglL/kn/LSl0AVHB6OSxn6f1s9XRHFoDuy
8evxW8GUK3iaECn+2CualTnW0/FY6J2HVuLdzyScnJHlrJ0w8hdsFYOJ7kUy+/v/uHUkQOCylhxZ
R9Ajq7xRN0dqxi2ufsh5q3Ybf+3nDJxiX4pZpRTZBJTstWLuo/lpQxUmEZ4oqy6cWhazuIWqNO+5
J2HpV76Ahp86mfQsCxd3hbGWksiIc8vln/3D4NbkBZbiti2vMYph26AFVma0RsnChz+hqjfda5bb
olkvksOGOZt1TsHKTITYTxhuyV5gyl9XlwP7f5Nx/sEEHWTc8o9pZ7IO5kAQYHuXtJfmjIMFr/Fz
xY5MHxk9tPsBa9b0t3Qf9y3aA9yVmlXoH5xOwb/NB3TQC6jMtfw4+NVY96peDm2rdCcrnnbVLTdg
ikcscI52nkdZYdt5DjcNzuHhrLU1z8jUqKXa9IJi5ruJtpOl960YCFk8S9Ck+hyfeJOzxRvSGxr/
+1vzlByw0Ck/eaxMIWMHQevVYdZgXz07XAaHT1uZ8817SFpVfj0qVlxk6Hc1XcZ+wzgLmLl2tba1
oMSg0EqKFe6j6zP4btR9ymmLNn+OIlCVJTi9FaKu2VuniRhUEdT2liqpjfnQFa5SVfEnrqw1G4k3
28TqjCyDIT7PPe+Oxysit+sVen6CDLGfauzLP1LHSKzWf9jaWLhsUbWCpSUBOglcxW3bF+fvvGVM
u+9DHfViKTWXHjM3IKVSV6DohH5g/5sca2rPUVw/kN1vDa2TSu6oK1J8WBrA1lHsovhd6Zr0J31Q
+1jhP0ArD46wYaBSttQPzvOApqiovf+9CMXSHx2H6bktpEWUB/Nvf26kO8eNYPFsMxoYkqOw3nwb
a+SWWAacv03s3Ba7VrBuZBxybmrAO0hFKx0iBwCZ6cxlz68VaMyWsXlSF7t08To+avcJVSvCEFnL
Smjz9rZFsYTvwm4yJuwKA6oZL0rBuXSl3v2SK0qSFECLgA50eGT473EZPxFMeeQ4buDAJqr84cRD
VK9Vi2mGxuEvrSNEo9U5flV7fHclVWb10TthJ0XJkehEzqplGM2JSeSucVIHd0u+C5T5bY+Vu5dE
BL7hqykoe67c+k9ECuT1yPh6e2yg7/iTpul1tD08tb/DYAp5mprxZ4AZhAhg21Pzvn4GU8gvKQXd
yGe56Yy3lgsAJjlpppHnJyqSYrWlEX11UegTPusnMJsSeB8peWkvra3bjdITIyNS+FpHteHXnnCe
LCUo7DiVMRzraGdmsyazBixnBSJSkIaa8nerZoCVa+YLm10veY7E6bJG355fij6vC7+4/iUZhj7a
Qog8AJ4b9E4iSeCg5g4GQu1L7q4fMdT2PH2X3OAAXa0fpQqs/RQ8bAMvE93RoGYEPLBi7hGbbeOg
mOBM+xxhEn/PSHRiI6bD4MxOXLUZO55q146tm5PCK8qMitw2CIOjGg7KC0KaQNv/6c5h0FAQQP5B
wpnsrWl2px44Z2D1UWll1QnqLcCsJax/z7W337g3YDPJvuXIw+nflAQk8Ni/97noxi1f9QMnmPCq
KpS8W9gx1160Qyw/tQCnVxP4Jns8Khyfn47ZyJrWJ4rCXuOTDx1eecuQqYSlGWdeno4rbngEoJbi
YlAUZnWu1DIiZTBRFx/6p/42iIVxe3nR4RczUgCj53TUE8tlIrIIWQEkgNhuT80nUeVkjdXGeGgr
KKFHOYVqYOaXMxcNkzv2++0cK3TadmCs0CG73we4Post9CbRy+EoDLiqUq0vgGAUU+0vBnMOZAPR
AD82DaX4zABrmwgtBewbuoEFyIBXdaf/uYY3q4wPAZj7yaWbGcizSJxVQRIrsGz5sT5sypZ4eQuC
piggqvIt3ShC5WDRafSYRZmeVj2crOGbeF7VHgr1wytXWPYVPXSTqrHG25rvcbomQna1fvgGVpk/
gKlYgADjsbV28/vh/zGM2t+N+uAdnPL0v2Z9pf6zbLTJezya1f9fPXZS2k/jT1p3nzjLm4ocG+7o
ujs+bmhpH0g22p64sM7pEeukT4/9N5bzbb/+8HDDf6trnrGPIMCcDnXMalsx3rpUKCGGJdUIvt/t
wDLw/IlCwLn/bjMKgnC1hfVAyM/73Y3Y1pjrfQcSigOOrFxFEzlOsI2r8xI2/InZU/2wYs35CRmd
rw7mAnOEjsLgOzKPvjXsifpuWJxErp1yv1rKKIxI/U6THN2Jnr8U31FV5chSiL1TsAgbf/kdJL4t
qbxh0LlrT+AeCNHUpfJCn9x35fGJRYVNDSJfoVxeYpTuGn0ExVDoWZpPn36LF83+y7VNQ2bGtE3Y
mH+5pePqwIxJX1b5XULrJCbH+72S2Zco1OeXfwyYlUxIQlxpQGPxq/mUndD49cfeq/sTfEE75tcn
ke0MTmPz6dzlvI/SEBgGkKtJw68YJ7YbLqEigzFK/2YIkbgkoIO+hol9ksLuTYZgBUBsulaqW8AC
078BtoWcnI38I5czG72rhQJ/hsVOIUOr/EqQFZ8a3YKd2aXNTTLTag6T1fA998hStAEZfYbpzp2H
wr+fT3ICfUzaePQBSgG21torSH0GCr9O0QxN+glPcrKSmu7MmSWJ3zFD18pHoQEScIW0JnCy31OI
VHVHlLGZTqxQztv+uFzR/SgGQny54CVbNflkRJ1Qs7hNHweiVgtqHlFFKklk39c2TLp1KRSXSqPQ
KoFumlFAaZSvRrwZlPBCd9yHe7cYhy/UnbyPuy6ZBVvNgsq1IBtayJzAzIAeoK8rpQeW6VVjw1CP
Wi0SdRp3dJR076z3d7YPqKPIZ5IHsCGSEr1MDZT9Nb1QxhykJCfHwReP9WzkYZqRvIB4lzSjlrcu
T+SR9Nq1h50XxRKy86h6WWPas83ili/uQVNRZk34QwhEy6i4wObpsql7Lcqr9MO6Sbl+X6SgehUK
YfYFTECD3agNXiztEW+bY4iwf5sOvzlUpSC0foaAOlMSO8FvEH7BdHBWr2xGArlE7qRGcrAe2IsO
8wYpMo/4dLxyrs2A4EmuNpKvP9kTJ7NRT9cAsWFg9l0s+QxFcMd+vh4kueao01bbczYE3E2+va6V
LlkT6f/lo2pHfHEktMavv2/DPdfS4lhDWN1G/u8iOHFPMta3YxIhhnysP4at83Fl/KXVL8rFOPSH
nVNmd4BT2di5i1JxwzuzJdvEw87dzgvAtk6kr2TnnONZLPOx49H92vtQFmE6jGGcBSWB+mhdymZ/
KMC1/0LiVq2M9p4Gq8yDO8Lv4IzBNj5eDkN9enHIGGzYQ/mjeEz4DEbedlhFu3OrQKyBD4eXFVZY
ME/fa+IDiFn6mA3Bj0rsCRBhcJwmfZYL8gvFPbPNb4UaCDq9hHQcjRuyUr+QAc5QLgPwQxTbIMev
IrSheaDpEt1dG7BVeunPp5rh8JrZndIeVtD7a/UpTGygLk4620q1W58zpYeBbw1gEJULsVZlt3O2
nTLDfqyDEJ6KQeN6pscaGTtrPKiXPOJgYcut0StZrjX3LA5C42MuQt5mt56NUfnsrBQwbJ9eInzT
/e3YZa8qgWOOgbOkD1XUDh38RWI9/RINprAiKAOoULisssnE+DL75f7Z4UMHADKbF0B4jtt74POA
xk9D5XEh+xNiVOufZzZfjBUkztw0wpJCX6iJPlelBVn4WxBzZwDYXAm6hHtwwdlGDBIEfrGPUG/h
Yy01r31inBVsTxMcubY62jH32Psx4t86bI1dBb5gOXRSflCri7epYzICZAFIaFBOzdiJpsC5ncOZ
khSoQ5AUFc4xUHeMJfsQL3kacE9L2vlehnwJ2HxwWu23ZMIMyEXWriPRWBQlvJx6ZLXzczvu84Oj
auM+v6HTsjqQxUSUp9efNqq74LOy3eunw261O0hJ9+WvjZZqj+m5C+TQPTSYxhv9EGIgH2iLnHUt
DPEl5LCpIhjpF7IWvdyqMUApTpnAATFkF+hAs2dMg8iwcpKJxuNAfNE7xdpg/fxXWyfMlcLszY52
BlA/x2bnEm0p5ff7OT0KdJh76NVZjuZ63CvdP7Y68sI2k5FFW7PCnyWajw40wtjkwt46Z0aAtj7z
8o+3Oby9ryB9OobLoLXQ4xQQWMKx9w8Rj4vbIYQRxjAZxJhZWZxvHnAGQsb07BSbahPI3Ms9l2rC
XJmT9LA/EvwYWBs08SSeliDiWCGYRskqa4ob2Rrxi3ZzKes8bN5gbM/Nkefxs8sO4GoDfxCre4Zv
Gu+2YOEDkUXbqVjmsi0oPwKBVL+H3ESo97RijDooj+99CNyqUpfbcyToIe7yYf2zKyduuYiidE6J
CWBTTFFt03XfQyIi52r8HavM0JfymqZEC5RuYkbpsxGah1jbVaYORYv0+mPlyoQwER0C+nBIigWO
R+BWMa/udjREU//q7FycHAg7KZT3aqLyjW5Kf7JW9q9ss21j2OG2gRF1Y7Kt5/56atn++DwPduZO
uGWzfIPMsSRaBr5C4X2JYSwARWf2QxOOJjePq1eSbotXsCmhT0A2K3rA9S++5ZWvZC0fpAwEkl1v
9xl2WcoF+IbMGA+gkOub1BtT8UKZMZQGF9niw0e3uSocibW8KMG1mIc6K+i/sGkYWN3OXKww0/6v
733EgR7T6MXJri+K0fpwOZbiZHEaLGE5P5Udj9wyrhs6Uag8qlkt2sNqwkwrDChVJR9QarWzG0Oe
td3pi14q6tZnHWukaOQ1Xyoi6J08aVKDejOfrWig7PxFF/2y9maKbQG/ifUAtYoJiLc4flfTG6UC
1VAsurKzzl3w1Y38y/XVHeebX7DKK/USlevJDkZtTE5MIBhL8Yq+7f6GDUmXpWZGD3CZLUqu6BH/
6EuSzahgYVzuNjmm7FNQNpCEZGyBjol5xW7mT4wQm3tneXMCUpiY9n+xhLvcbyMuwhiYdFKXSAyJ
ivypyfnDVQKarI9OKXLRe+274rqINfvTeoWRy8i3YLriVa2a3eQzm2ttU15+yTH10NEm4dZgvb0b
jCG9MY0LgxFsTTjPr31Sioj0vF7Fzpa0p2tyTslmJvKBlFJADp4X/P0B2N5tOKfSLj2pPjDop5LZ
uxoO1wFvu/NkxX1gK9SNV2fTNPcs1LMpoj3OR2oM4Heul6N7lotG/K/IzEiTfDKWNnHblpveYeLN
Gns6ycGnDixo7lrLZS1gOZT0v8OT0uOCBapPbi68b73ecOrzR+SnwhmFNINHPRR2IhIjk2VzZJPt
7nh8cUEvHB4bf/2MrSVEtTXbTlFFB1UzMy4ZkrgLISjbO4KJ5XpQL6N80mVXb5nSZ7NnmhheX691
eDFC2NC/o9ho303f/gBDU6ZUKgye0zSxlvzS+jyaj9tHpsERVi/SUI1WvXKTODm7lW/TnwLdEGb0
Fu5zLcKgLWXTSpvKZN63I+xq6cLA0IokrgCzrxIyLWvzW2EDTtSEAxtnZ8dK9Lrfm+ALIRFcmqC3
jWtb4R+RQhhMqE/Xd4hCTJE1PzsM0McIgRu1uqs51qSxqGjezTY0Sa5qi+yZcgBolAUVKgBY5cok
1mYM2YPUWtXzublgo6tymXXoEtJqG9ctJYH3yr/2s6Aunqrspawsq6e9vTiuZfleRbc5eMjkYPpE
CMpUnlT2OcZ32UqDZutsbf1cAgX0WkKWdUw5RobV//ma/Qn7hntgYgH+++nsEfoaMTiTTmpy7CCF
2shQA6LvSrDf2QyBVdyf1VGUzFhiXyqJ2wwddeQC7ZCcaWhFkXtPy+lfEvU5QlHwK2NCaVl1Xxv3
EnwhvCb5nfqQJSsr0PPLYhCRlMOEPfVPWLZW+339ZCrAcL8/nV5CZVFuPrAX+xGa2b6H9EX0RTwo
zWzSo7Z32qVCeQgSCvdHt0QwMLhdtdWCxxCD+2aHk3llwtgsFFhC073oCchaUvgR1sVeL1npf8t5
STXFebQae7sv8QH9petAqkSk7PcxTQUBrjHC400CTuTORF3HzMcC+abXND9/WgK6wEhXSyv1VqWE
0L6byb0+wUDfR/5GZgviWG+kyBpjni3Rjkz5rs+zDtTKnYSnFVhFTTI7HBptxsauiWMcYEHg/B6g
yvvqVE+KePhXbvQI501REBGsUsbCWBPaSw35HTp1zYFQMDxm65PB6kkuB7Sa+R947u5kn1FYVrte
u55f95M7k0cscHFNk4U+1HRQFHwFjq8iAj+zC7dqTrP2PPqu3aPZPsAfQCJ+UnqhhtaRy/MbpARq
nq4Hja8eQPlYGNZX3il9NB1eIc5ZzyOGRAGdJc8qlKEfBt5WJLxXUyoeRxVoVm+eo8I7ApRDyNWt
msf9dhaDTilvHQKH75fdB0DRQLZw4FPTdlM1E7jS6NjyNMixPrI2WB2scS+g7EpBGsTUigMKDc6H
q7cuvqfktfpSpulCYK6R5cOgTV//Lq62PfuWtqZrKYA/qleeGXI8NkGGXaOU/jiqFIloyhGfdwGa
DY+5TU9MIsJrkhpW0w+DwQf745MuY/8eRxrocb5k+52ttDsf/AOGv7xdezjH+vcD+cdZQEzbzWsM
Kr3BkFFEFX3IMUMC/f7WZIKPHEGdHiNlSp5Z9Q+HqrDOs5QSrQ1Hkzu2i5T/2GAzZSaw1aoI87vE
7eqX1Nu3IHTYAJsveSy1HI0LH8gN3tHkLWUvKmTek4sIXX2YsW3eel8Nvp6bZpxWb+o9VTRqzNhV
YNqybtj40oFt4bapB1FOaqJI8+SEjW+dcbJYIWYvsrI+YzKOEOdv1qo4rXRBIDrp6ZrVbpwvBUvp
N9fNpBMXGTAnB5cEWzAQxszVPCFkCRQzG088BcCJKY0WQbPRD/jC8mI0Jpk/XAdXTSXSogZVEJuD
1FCI2ikDtpogutbORnPkEKKH5C6N942VlfJjUNAUM9UqaIu46K7y0kjESJvTYRCu6iEA7Ickkwot
zifw0YScv28p6OleRjBPFSDllcZjNUKRfeIQBakeGnC58IlS1vQJTBrrCPxFPcGJpTJVUYb6w2cy
F3WRh7QphKT3WAnEUDJDguEohdWlmUZ7TmEiOfx0I1Q5YjHwVAT+mOpVa6MsgeZtpsObLu+O8hWN
jTvcIfbxon3Atp0xVN7tYCpQalmRYTlPv8o8YG9At3wCkcz0NfSZHRRpZ+MG6kfkCsfO9lh0mlzA
iePiMRkArbJSiBlaELvVLVi/gI2qXCgMu+KSkcsxO1IP0mCuVsWS/A8ZtdhSEwJBFTtFdP6iqpiK
hitbtDLd2Db0iWwQ6DSu/jerPpFPUqASIVyAv3oqY8rvvTPjOhC08xm9z0w3F6Cr3Tss4SPzJnKe
FHT9APT3t7itf5L6GfA8ER6aLQmIiFe5f8BjICbZsLrgaNAftjMDgTUmyTZu2DflZKIm9QPUO/PS
7iVyASM3yWVE7a4/+X4pLagt+TdwbCXLmgu5f/75y2VyYl/mdht6k5YF3nxD9Ty+doc1y2PfSNdJ
btQZHhu6bULg4qamswS+H/zeT1B7RvZ7Hmn0payTcyUKvBQC/eXz2RPe+Y1jhLwkefkxwjxJRRPy
oFYhNhp3wn+1wTJ9Q+Eha+ee90uz2Rn6ZFsWDs/iJRTmOWhMqZ+HnwHuqBFU4age7fj/dSDk+JU/
mYzOeuYOEt3D5MQkysBgfQJEj6hbrm9vf+js56zjR8by186EnJbN/clzASYJo5aZZXzi+EBuYoWp
ItRH0eU/XcuPODHi6afzTqSiX/6chmtoHwlsi4EvOBfSEMYVNDtNlcG1Fzc7povuzXqSb0lQIxOc
7sjtZJrZEwRrTpSn5COVTqEj3Bm248mY6XfexwT/Sa6SC20Oa5h4Z8pEFvT3o+i99PiCM1RY1aLz
nU0WGXvZdeKHAZKPbekBfCJCE0gTr5/J5DOkAfIT78FLxCqu3rpAhckxo+VYkUdj6nq+412Uc0WY
ONDqa2/0mQ8qUw1SHlxYVWpJmRPsahoO/6FVTWjnU/o1XQ3mEysJ1WSkh7SLzyw5V+Y8RssuNk0L
1WsLcxuAIoxlR7tjSlRAAo2SeSCLWaI8NkaPaUcrE/pCfl8ejjGPrOI4NwmbRi1sd7m7ng6Ft6nq
ehtPWbT4hXTOxn9sylY5H4j5Q1SV1+0hIxcASwhK+L9f4ZhwHxi9BEaNKzsGIsCgQwYpb2UY3aiE
S5M4SNmx6KWFIrQXihhpQmdf8JUnRV9jUBE5Ojo8nzCYMC4e5i1nbtjApwE13LfIL+V2xkT57HpI
c4mRemprgLz/u3xYlEWp1SB2jkbAnmZkEvLwJFGEFYwlZ/DHZ6s9uxsz6bPqFG5FIdvKtPRrOmIX
tFy0wKLyW4kqvJAmFavryvwmcOVkvT3fj2pu1oYMBVPMFsxfft66U+LKNqpuviC2LH3fCY5LS76P
yMOJXz8kTp8nf6Moe9ZYNJAKbrd2uT0AU/K0c3AvItw58w/cYEs/NH4rdO0LTzUBQcW4oGEn+Gm4
R2PpMwzNBekrFqGQAGfesXCpnEEjvT2UYOua4G2Yvt/W4Y3RjVCcU8HLvyvwUdl2QspXbxgJgYol
8zZXbTinSV7ZTWCVCzU9gXJtm/g3aXRRkNUsNy5fNEJMn6OmDDPydXsnCaZBAmaY2+2P2ZW2yhep
qEb9ZKOy7vxI5QOA76jR7GvrP5cIpx1QHl/aePPaWLeWjmP9n7ZZvLRXQ2Kr6tmNGG/7Y57e9cQy
BE7UL03uYNdo9ZMvuyAw07YaJydjUoLspjdQC4wHnMsmsaoAU0BZ1/NLexx+EdLkVLISYD+UQdyF
1Zvt31pdIzGbYMZidNkdjdLD8J7inTbdoL/OOHzhscuzmTPTQYWff+Hze7oyGeyLpmt7/GsQmDpd
9OhsD/IRSg1g0yvz4kZ2h5bcwA2CqZJXkeXRRL+etJRbR6P4JiGmg0SquCk6Ov0tPD0LKAKA9FH7
OiWAsl8fQoA2QZgxrZ8IrnpL7sYpCzy8cC4Gz89tbzpavMVjsDWbO6V1fKfNDSz61JJxPdIGfyBH
zcGZS25pgdaxAAYLRe8n96+sZbSaGEwtoZp28czfaBkp+0sTBolZ05xnRENyuyd1QMdsl/6y+VFT
8o4FHi0GhD1LxwqEE3iTQqW2el5L7VjBKvIByc18YOe6++wSwcXTdsY2oNu6EC6wPRb4IR9cdloU
mqVQT7IPwX+bNarNMhRJE7HhpR64E1tiYcUym89phhzSiEW2AzGnEc0qyDnMMRkYBR8LFH/24nK4
DOPVrGP7TXIwDDyAVoZgGi5H02cEGbx2GF7QEa4do1jcez9+/34HzayzLs2G0shbdLb7PV3V2xOq
hzN8/AwvGn/iU2pGtAWAIjx5zqv7eT3vqNLYe6hxkDMP0NPvrHj0bVBdU12KXWYK0EE1VAKx/FVt
pNqskK18EZoFU/vK6+5NPPMshHaL9/J9uuEYk73l1DGSVUW8dByegC3ThiogVkliO+RfFx4K8+mN
kvljkXexGMqbYr7K9cp123J1kmxPxiE/g0qnkMbM8ivXpgB58IlPQszZdabnSK+f/embKxpVdYBw
F9e8onLW9JljZ7eRhxmsVZZ/x3uAE+hL66FcDVVeaWAM7isxoT222pZl/5ukQOPW0RdugCUIN4Ad
TVDolTNLaJJGCRVHDeBVBDoAl/2t3mTli2Nw+YyHhL6+UrlgvjQp7EhdS3zgw23LK821UOL09af6
J1ZVBalD0cfPsexdKpZCxRcIfjtiIKcrJbwtDCIxF97hIDs7pIaV07Z6AVITsEfyJzuMCeGNyKvS
yzPOXCK8o3qT3F1ZHH0U9op2eCLGVm/1ZtA8aeKZixyOKcQp8a0lLUIScG9OnyStlbCLIFYm4ToQ
qUUExWr6a+aALeB/M63Rga4MAwdDO+K6IX5KC+MJwJKQFhWONt96VuYx57RK3ILnt3nZk9CBFTaA
rP9d62nqrzIkXYEFF+eTYpOQTqNvf9S3RbsULIr/gR9aiauwAGA+lWZ2F8npFjG4V2Fp4xH1y4OK
D6kvsmagLaHx9LGwIPxoeU2tCA7IwbhOZ5JJBxOVpUDOdjSmPo1E6j3aHUxmGkjOKoQhn+336k9G
ZyCe52nr7t/5Ic4NSBshHcLEvPYxd//cBaN/d7Cg5Ol2SYd1KOEicdLSuZSVpU476uGw6lGpF36t
z0fC/bn6y7CX6B8eKL9Xx0AoG+VLp2b2phRm4jD5D2q6UxGuz/T3p3xE4DPn9S+Hd72pjRRrqk+l
Io/bWUjYK7xIwwrKFVP7/6DZuSWY6GHY/tWlRE9FNzaYLxkNq10PG7cBOHF85mPxzZeOfb+45fsT
cwHxdA61h4ORI2iyBeK8kYBCTft4YtMgiKKNmNxcq7Utba6OHyJiNDMdEh9u8Uw6RH5+pEk0pE5f
6ChtwyRaV/dz0Bw7eUCsugg/KqTPP+4Z/c6dvkVO+zU4Doi3dzswfZWiJmgndFzVsGLAWnHTre4X
kW/ONNxJGHcORHC3Fs6QzaNYSFDQHg8IQ2HSQXLxT30DRtv7LWE9WnuC6LezD4AT0i1uTJBMUaHf
3dExWq+2zwZiNdPqnf/fJvcpyW1kwJdu9U9PfHLewMZ7Bb+eWGZEKmSpuTtHpikxnSykNL/cR2DR
zIpZa6C0qLJ+zmOSDhq8dl68xzH6OIb2YPKcQh+YhiauEGiAX5FgVmK+2AW2vA7zW2BYBIozT0oz
UmHLLIL3Ts9yqCMjOQyu01HFnKbROQb5rqflOmm+Le0dQMzfWTOrJ+zYP05rtDBzz103O6mKZ4XE
AMkn48Y/04ZBV2JpSGeSDYXozjuLdB3iyf8pwRLfi3lZ5De4FC1eLMsSRJHT63sRcnlgDJoxwnaE
tdL/NbGLoOqrRMrUdQdUPOmGl1duoCQj3loXOEw1Fa2rryydSjAjjT/WS1DX8S4hMNqiJBU9dIFY
D/b3pkOzEJNzpQy7knuxoCzmHVJot1Hcyepf1sUl2BSJcpVNFXiI6QisSCrf/1pLm+bFP1jjQQqe
Gx8JVOwOqtcySTnK2UYSTkGep07fcUXABpi87fyTDh1edhcv3t/Eof6B5lcjDPTar4i3w0zD7MFX
wfPNdS5NzMTZtOlfAqyfEIrniz79EP1TARGwFLGikx7wWFEfxZqmhPe3vk9CPE3q3ty1gEEc7DMm
/Gk9ZNdg1TGXzoEQW/7mZp1PQBTFAKvUPXcK0vvBgyQ5g1IFJBhqPnysbEYuqF1S8X8FsXdQG1mW
m8HO8a2YUu2NseM8QcjWGp3xK+ds8OJc6LeMgfIdP6+9wdylgvAglLkMHYvnXVz5oxkZCPJOsgw3
tuhGZawR8y+O8bhjbQS5ZjADQ13NzmsGOpL6c9gVUy2RBCbvlFi4L8pbDjugXbdfCIQCSYkq9zRA
Nhn/5SwunmitnAK1a4faiwHwtJFnrZcdlcPlMj5ZEIYtE0Hjxr1FPPT9GidVZ1T4FrgxYmUmt2NI
JTTRRB3UDKWxyOG4/m8/3GIukVG0IkwDhHPXc1D3jtyECCDTchxSTsUEAtwEsokFKYIP904M8ZkA
PglMv8CZJFs+YoSm1gn3sdQjOapZqdkM+QB1ULXahBjT9QcIjXbKnht+r2DEZDp4AHsD20oMo85U
OtBX7koQYvRIReMdCqKI1tTdtLB77X4cpFHhc3c5zVvfMpKb+DlCwr+/eNG1GgvDUiWhB9PxdhCF
0jvKdGyBZnh3+JE3DX1Yx507Px3qil/KcEQoqxdBNRjYw4Q7WIckQxGYdaNjT6IFxmEc+Vsjvszn
hBPqOXufeCmceVezfZWk8U/0H1uUuWp9EsYUSeo/Pz7/kqq779CSvUwcPXXPFr7IM4aDR2cO8GiF
C8UI5YNG4jyTzMmYnxoEXGQCANSD18mZR32u0dFld/MxQ0xcdlLOQcUv9/dbZ5iHqSs7ErHFBlF4
Y+qT4HLp4SMm0ZoBEp7essAsmQZEDI9XnDpu60/wPpQabxFviVwycG7e4kR83z4i5OjCvDHlTCcV
bxFtGt6mkO223eQQNQEUTRc/yOUstZUXhQb95c5COcjMI8uFlrZyXWD/LGo7syrqZWeX0lPU2lvF
PPiEtFPDoHGaPSZUwOLParx5mtEZY/6Q3RIRg/ru/EhYwL4QBWVhj32ZSyj1hKqGTw1+osAUK+6o
yh4Y4vZ6/l/aohe+NwJoSLzU2flK8L4uF4JLzl9/xgtF7O46xJBOt4Xeh367782Y7kyF7TzMZIvU
ZqZDrpldRQESpjGOk6Gml0zV+c+b61Z0OKpuMJBu7KAmn7SP6GJ36ID3zlQV28rU1f8hemr3JeP5
Kqgpv4ibtCUme2BXwY7F+BPfNA26Yms8zWMX7GV0LyIxv8qVvtIrJI8IyrnTiQreBwJMz4ha8XF4
VZyuMlYVhbK5UUC73uqeWdpgbld2YajMq3vislEH/WUI7TnHpWckBi9MjlkJXua5xPGrBTzHPSEj
qqLyzpaD06elNvw+pZ4yqo0mzqhHIeGPAyi0Mzo09O6dJNPe8UPmBwNNgcMBhY4P3UgkJLo5sPFv
0eVAlFLx0OSFO2IsedOH8SQPRcVlSYLKwYBMTflDkXeLJsR7seX/OkWL5X6E3AbWf+B+FWV7nO61
uREwtTTmvRvvSjG5xN/4Z8+utP9lEmZrUhIM1mPZRONHH67fTVTQW/jmyqI7qq28fSS7pVGM3l6d
G38+tvBD76lucHxy2HnVTaIIynsPZIHgpwQbC7EhaTVJ0YQKRoorgUFRQIMYGYU4qdPKiVpvhaCk
GKqGw2qxqlG4fYa5QIM7EBOi/G6ph0tgNBbdyRXPnCUarh9hx3wZpBPLdLGwcQUIyNnnHLRJS9QJ
NlQfFifjuXhvG5+9KPIr/zHVCxlxRISq43cyV9uT2YLr84ImnP1KWIuwVTA01Sr28MpDVSVCfqK8
5IrA1ZqI7RhUVoPYJuH3xvOrJsb7vUjveWRz3ocInAvX4JFkLsqgu+KlGCeVvhsdoa+6oa7yIUqh
KgkL/7kGOb6rcdcuNA3HHv9zpNgqqT6ZmSXOiqi431xMvWekB6Nr2IwyEmN0W+hwZhNiSinOnDAL
ImAwZBGJooXjPRfN0Acgvx+6lrR6qMWdZBrMarK2UXvWWrt1FjVaakjl8Pif7U22959ZgVGUhMng
D4rJT7MSvOcc80D+e3OpXHR/SlKfxfeXPJeZfjU7DeDMW7GFEtF6gfB7qg+KHpZvlTcqDGdjb8ia
bdjwQWMqp1yF2VIrBVIcP9nK/AxbHrNXxfGM20FJhSFx09cEnZNJ8NNB3+mBRZnV1E/pH2T/bgz4
fAMMKN0IOfuWiAH3L4Pj/6v5pHd8BKBhAk2poLWLODezstQZLez1Ys9lSzTl1ORrkOYzRp4BFdQ9
lYBjmGF6xMZfHbtl/p1S0dj53YcR4cttqszl47srj4+FLST0ppUotu83HIUPw8m+rMhP6PXlG2r6
mAyVYA3i/Hcu+DodM1YmELctc5zx5/BNawxLtHNixUrrCMu55IIDzsCrFHTRYc5ngy38J3VgnXCZ
eEWirn6lP1lwZh5cMVxM/Wv+wlTw1BHzxjU8PZZms1L91QNCak9egNaK1CFd096O4A3TZHJYH47H
W3Pl64qJC32uXQNAqMKxi0gFaTHoaCXpbq3Acb35Pf7E5mKG55ushU/uAm1ygmJxN3yO33BD05vJ
cxZmo6j6QV6wwzmeJZkVAjuiCft1ka0NPdh1hKPveVtNniEd/iFaxBeyj7u1v0rbyAlvkvZneiLW
/iCsNTbTG/mAGqt7MZdZxRnYGKFwSvAQn7pa3rRw1e/MpkCsIoOnBPuoP1K+WPw9awATvQOckEbN
kL1y76EYHtFDUoN3KeRg5pV8tbVVz6T/s53shjib8tS82+LO9UpAdLMS5Lhxob6prdhQP4RwKIkQ
51xGwiovhzy+nyDKalwXnL6CEheKrykiGFFSMJWlQo/sa3Yc/eqwoJ6IZGasQEFf7eutwxqlJbU0
BbM8LN0he8fq6ktGURhhEUmSuZ4Hod4e5wOE5j+q/NggeWdI7zFfI5WJwMZBiT2Qvd1w0yppjwcQ
e9nhYwaRyAzXioVjXaNsbUl/cJANQIsPwFhZQw8Vbq7PPWvaSlL6uWKYshIItC6OUOFL7BdIPG6e
E36cAkzQE9pObWZUNrbJN8j9QbhhfPiM3DQdBGI1SShMynvUF7Y78s4mduw/EZF2XyhuZROVIueU
AwpVaP0rE7TCpFhBT+WAhUoN/bqgWX4ZATQBC4Jgf7yXadO8JxDM5Tw/DkWlp2pkMYcy3+QgK8OO
CKOuTCsW4Lvo+idB8ImsYtXqqPQs1wpi4OmABAxuqFQheT35POfpmuQfmIHN16CifeUR+NwDEupa
/MIDikZHHk2uaoHqcRWcdTOtvjRkwJblr/YCSGV3wLnl+6QF8PZNS2c4E2Te0OWj2eMJJVDtMbLk
T+YirOb64Tzrv59rRDpt0GGppuJkQJwpvOI8Lj2GHLEs2tQzrNapahAaEtaEzI03CfXD1sn2vKro
RVMybVqYL1315hrRpAvc8hfvGfvMp52Ka8/Rn/AlKDiT9/ifI1/j/M1/8+f8yBFoyVku7bYv8CAI
ZJELpArOfRhWc/oiaVY9anSkmQr2r/DgZwow7waE2twxKWbq1KaPU1A8Z3TJrpOYTmAbVN5vT1fz
r4FzJp6G18sAMdcbPt7+mGGUa5adyciPJu3ElrpT5tv8pNXHU/PDuuKjLq/EmyOKybpPFPt893JO
dcBU6irhViyjGbEmiS09jbYaF0Eiz9mi9jmiMYubyV8Udz7rXqX7/W0OVLbRHBft55vg0sFTADV/
vlfYXJ41JUwMhDSfbYcFiWAQ6KlvpIgbfgyEhg29jbswpEb8EJlZ3TyLrelhCykpw4mczDBw6XI9
q2VGHcQ5E18tb4JP6y8obkAYGo0J2zPKUFQ4EiBZHngJ4LFA1H3SKmq7/0zcRWscvz9ZZfP4i5/Y
aBVT0NxiBK9UlAXLwt27nmrkjnrRcOYkwmHaKl9P1k3DKfmd6cXIs3eH2OFh5ZzM31Jdf9GPmYyo
VmG3KOdqSEkBEWKtoB/GvDA8t44gsQ1NeVQr/eDoNVYlTQ9x95zaaPeXabYWgZds8aZmonhA7JWP
FGORu8q7a1rYib3kn5HEOq5rtv/MH+VTHQkxErPwzihDq40+9BzhLXM3Oh9QO0wW9vk5xG468WRV
sStPouNfmEwEw8cZmCIEBojl5IJJlmEOXOYeQHgEPU/fNukCB8vRxvH3wOZBMoULCHptYekFJvGf
HooHWunpiHPgrbmMoTMeWJbn4IoSBjQJs602sm0M7cUlxzRNTrwy+0i7w5uji1rn7FnSnOjdfg8g
DcrsSbyFkPqLDzzp+SFHM1nSDNAqVSpcD1G8oZDkyJgC+EO9iHlfzhDNC8oO0MHk0ByAL1LOJoS0
bVbuAkagXBFPmqqzFWsW0S9Jyzsf6cmiEzV/3yPT8Oz7psDxvjMRRgbRLxxVHKX+pujXjK/dWS1G
0Qd7+YsObwsg5Du3Pxvg7r3J45TBnh/t/ffltFX5VMLEZHFj/zk181yVeHGVkIh85O87nm4HB0v7
E1cHzOF5XFz0nfIOhziJ6cOyplhsTTZkrAu3qpH2kYwFMiwn74+FuyXI2tg1jtefOZyZOC3V/GGN
JzItVRUSkZutUpCW1/BPzcDAIbWegY2ccXFYB8pAxuwAbVXxnF1yArvGTIh33JfFhniYPi9YDoXk
tpYwS4DNyHBaOQwZALcbLrEqzjNKMBDWsB7kVrtaDjs7yGWZdnE0kOM16lV0riKGZjcHYsaOHXgJ
mraqStS2vjADJ83jtxmbqePENAxTOwET7lnTJqGRwxXXtNiIFPSeN5TgOpfuzCD3J+47omtyxJAd
F2OIrzJBI0XaYcRqaT6+44uz43D0O43XQ2gl6mT7T1Iiv0aku5/UZ8RLW9Lavn2vtbb6OdcMfqnT
Jb1yjWVgxuQXpKOF9wWF11U5QK5Wr2MeXjkOaduC0LDySJOJKBbq5bc1/QH6HUVb6rnkpj8bwpp1
59A8/uQ9CuaUAaNHgXdW43jiRgu/MNUcSqk7CNH3oq3ESy/ZXGwypI6DGLsKRAZMcyRsmNXLxpKn
yeCxqG4MJUYfufgtwGXy7MskNkQI2xiYtp2/k2fS6iA/C+xgawBrPYE9/QvQ9hoTcCcCrhP+J/Pi
3+2ppWoIrtxHQ/t+F6z1/mpDCa1E4/hM6MhpbbibughzvQm4W/LdhQmtOQxumpzpAwFWugPjKOPA
K0VHzTsY/JDCkcWHPaXtChsmokY0QAwPig9pFkv7molx0n9yWnKRBUouafpYAs966BTIFAshGmGT
8xnE6ntHGCJ6iDWsOWsufNPH5hQ4K0PjAmy22Z9xylo0Mri693/u6RHW2xydb9CElTaI7XN6cZEF
Ey3EukrWOagbC487btal869Xt+hjVpL1qtjCKopy2p0GPZTzaFGwQh/Qaz5oShUw4dx7sOO+9Gh1
uj84HilmWymfLV7o787pVH4PKqYaPq4z9RgJo56xqZjK49WR1ENdHdFQDBUCDasL1oeTzdnWSNlH
NxiATd6EstkgdakN7EpnNOaYVbekKW7ahB15sG7ZdBwBE+0o8xn4pvUB26zyhtOkEKBXMZZv/6YW
8qrXVjjh0kuGXyy4AnTZB9wxKPnF9utrUubUZLoCa8QjtIK0xCOFuewYPDASq3P1kipSS8WrmuDw
YqvddXmxoloIZJ8B1iOf60xzOJ/EUSZpFXvjByOeKBO3RHEYel5C+fTg45QG3osZiqhbhkOg6SlO
FRqPggYrwwhRkBjRjYYsnCd/g2gfiwxyJAXYTZ0i+XIB5aaGEP9S5LOk1WGAeQPjmhtGKKcZgXvn
aGAfHXuFiTz2/B3XGbY234vRtMnAVxTeNL6oIlF5dsgY+b20wzbhmhN4A9L8hcDFpyMEbinHIoxQ
lrzbQx5vHA9ldD8e176zB+LfWg3VtlLbH1WVGnbs9L/UC0RxeF1exbjrKmtSKC6Iw7t3q1z949Fd
CknI2H20Js6xt9oDJ/7WXMgtLk4IUGY4uTDkXB7Kz/Fski8qfiKjP1azOPQBv7r4VRnXBK9Sqvdp
QOfMxiT5T9Xf1NF3BYne7J7UKBPIWevTDH2Ih046y1GUdsyVyoLZ33Dv/Q3HS/Ywtz6jl7FvhPYo
wMwydxZyz9qEXJyHCv3ynABt4IKYOvgjoZH4j92CCTapEYX+LItRaNMAxi7Ike1NY9hP38uZtowB
+LtAr1ikyag7O6r8v4KolZsDZBRlWFZYq0Q+KxLPWz2n5IPbt20v+ITsu5nW51qWRfp8hDaygk4x
v2XzCsq1pBCFFUFPKApAbm9vKCE9lHS0d0K99hM1g//MQCkRlOOJPPcSKSmfwWILWzUsWinmJ5Ku
HV8nWLQMqj1NqGR7MNyw/dHHHLCV+T4jno1CYeM3XouB9bXfi8f4W/9hluxq3Gi2M+rgx0BzZo96
u/MOidakKrFalQhRZf0fupxBQIn7ZiFbS0A+u/+7e4EkdeSp20qush+3+kfOXDZV02Foogx2j0DB
6DPfKXXVFVsDBFKHG2X7QrtOmSUTxvAbJciO508ekcSTY9WGnlBNluHvaYuIBx5nPUd1f8MuzGhi
R1ZES9aqAiXwekZPEeP7ByWbG1JQNQUJTT7kuEDRLrtEqAi0vIGNQabFXgzDhQ99rDE60VsXv1WA
ey3H75LgxsZUMc1nsd45NxjO7AWEYRWA/wrJh7um101ACAPmoRlHd2T4iiHDOohwJ9buCpVMAkr0
Jf3VLRVpIA53kEh2Swxl2hd/yhkozfDzMNKmTAkpeHhzsOjdrt1Ltm+JTfGAUdb3a1ndv4GChxDV
fX3wG/ljZjYZvgCASoHQdbkahstgljdsbR1XIlxGYqZtzE8Zeg/kD07Peng6gw3pZp6JzDnqhu0o
23Rg3dPrlNhl0Bbc+VzHweYKY7Loy9irr7K/hoAAd8C7PUXnOZ5ng2KNGKBw3tpGZ/lPjwiSZI3O
R2ADJR00GLUNBtiozluRBSkpVO4qzbUi4Qnxt3vvUIxeDUANb/WZ5noZO4AenUnl2F2KXb/D9Gzu
bQEtJ7XB9eW3fzY1gCIlTjE60ylYg4onDjjktaXXASQk9ZtkZ5kowz80bh5fXQe43TmMXCN8mwT3
/dWLDZodvETKJOk2iu8jV2/HhrK95ojkqVJ3TfAAtzL6MQgSnEk1We5OMZy3AOXg10rz8tzbrKtK
y/zKaCKDNY4VeWO6or6BlprxcDjBD0cE9PlOjC/Vq13zjfO6RiST1iDRBUaxalflOJ9eh+sMVUvx
/aUWvEAN0aM04I6uimtRMXm4g9LAzXV/OSWUNhUlOIafvIuyyN82HzprcP9Qs0pJIOlV+6zGKE1t
PFnmCok/XyUxHkzYvXrYZE8kJkVe7J203LWol8XRVZg5XavgcFTR0PA5AQ1e/7IwLv5I1IS4cTXX
yZC3BiH9daw15z+MYMIcJTK/ASC++tOotl/wPbuHiIQivfFYM0JpwdmcigXWwawCJIZ1hjAhpKRV
xoruIpbstNt4NhQKXM+6h2WnJbBpdsivso2HOHwzgWgwQYa1aySiLAZ7GESY7r6NnElLRdHphnBE
DEjMogcrizmTFyRULOYS2vxRLYqNA0oT7+cvz4xkkQjBfT9exaUSlPwnzQGy9L7Xq15E5hrTTCy2
bzITB1fJeoOOiW2ay4pPnepAzhP+8S+w+QNNr/+9RcqiP+Xfh52ycqeTl3IgeQnF3TcNgCWcjQKa
egLVRjqoZjfdRZ1UxhUtL9ivsEvYK/g5Uo4alcTBgWdGkdK6A9df2DcdA0lJXc1mww2sEDzI96mL
ZMBZmbDfZ7AQgxhw9yfQfD9JCcnMKt4xZVUenPpKC8vb9zBFVt8ATgSqpM1p/FkhnhyP3fvWktRW
zLKjqLR1uSThxV/XOkqUgSCHRboult9td0iybGw9FUUtc+PV5pEpLp+sOiV6sJ5k2NjLMVmQO0DJ
sHeCNEjeK0/wBY45xdnQ+ctvFmvZdWyXsVssuE4za6c8bw+119vWvnyE4XVYhvY0K0PHLQSFYXkP
nL5bjjXmT1WjhBGP2zoHT7mLSxq0Hcnf8v1+OBsCci/NMYNLiHCn4dHqUUGIOWgc03WzrRKJbHSL
eV87Sm4/nBu/7Z69xOAZZEn6w0tdMPhACox9izAC0hlQiNqov5EOgRch1HA7F4R+LRn3IWxhS6sg
M8qGszOeCQ3vno8HvfANfgLbu+dLePcUp3ywO10qIYrX1Q7bzqzKnDAkTDccDRWjqqeYM1ZI1Irz
5CzFlw8bw2xTQtP7mP9DUvsyoRPReLUK3ouG05b4IVPMiRK1cA2l2Uv25E5ktxARX4MV1aeDCmT3
dUqKEHttaK0QpF2rh/30OqxxKkD37+p8l5JGHTPk7jNRgHMT7S3/7R7d3bCkQ3IK1hZOFyLQC9dr
4bSP82//pFnyc9KjRxAxGsbn1JJtY6lpPL2lE5kqlAvT60n+ViY+0FMdddeiznaJVxhCzJlScHT6
q3h7nBlDhoY7pxRvknezOTYqAY5UMKPAmZS4EgGSS8Pwt7OSqdVerW5NCjcUTTznJPiYEXJ7iQ3U
DRCisO2PiOtuJTr1lGr5D8jGT6uKSoK/y6S3hl0WIbum57ZXiyoKC7lZZXZ8P85mvd4ez8l5rrxw
5ovSCpDrjx+Ut1QqjaICxEf6/A/eRZIkD6MjZrlzYE/A9FkRPANcJJ1Htjj8GMpXHuKEihxMBdH4
86AJwbw92DBLSNtMnZVpSUUMc/B2MLFRWcYz8lkE/UeEyzxhSTuKKjoBGIqbO7c0RXFNkQUeZptJ
a4+c5jhb36mM6OYD2eKPl+9rv4m2e4T7kRwKlkA6qmreJXkIHZ+hW4iHO2jmaA4VfOPeH2DpwoGg
PI3VoPVnVVfql+xHeRhsvTlBEPBDGh1Zk5s95LyBI9IPAMROvai+D5fce9+td0jSwtAGwbgHgefK
dB73CCcgUiIzgO6OnlYC26ZAE/t5YT5RnVuzOZkzY9jwz5Ryh/P8G/vHJUyz8EatNCz/x+GfO5/8
e91iyfIBGkq7KPgJum2VsgdLHw7EB+6X1IQW3PtumgzogN5qvDEdJiftBxvexqiNucJXipEJafLj
TXZCuBn3dgd+9Aw20BL8zqjGgEd9oovafRjC2D9KPpTZ39DOs2WCI5WAAdiAMwGpilYCz4O9pRoW
NiY8fUAGRfcyBeOxQDZYbr0apw5m37yN/gww8zCCxWqhMbGv6TIM5SW7h9JnFmmOelrKWCOrRBba
zNFC2hrF/+57fAzV/h6eEuCoorljD2hpx2kPhmrFdat4jCnGJGttSfyNO3grJaJgTMz+phXixB8K
dUlEHhvZm9IKDBgmm2zKD+v5+ZlSXReLeaM6/KQDeQke59zXv6oWDuGB/Kivam7uPhQnb5HgBgfp
3d9YBjPDbknZDliuuqUlDrpzEQzImkvDZa3cdMa9fGW0PjUe2C5px5iqT6DPj/R4ZrE6bj9WvJpg
HMJ7hfCJ5DOMo8Z92yODsSejjMHvs0i7BTOZ0t45CQtUIZRlKWe97fsI9leF51/n8Gy6jMFkMtBi
+IEu6OZ2a2eK+7qchm9lwiZFxjTs+Q1lq2NHzBw5DICXRyB20xOE2iik08Cv38KhRfCRFRWNl8qM
XKywMTabL85AJpm0g6G4h9Wi9W8rScHHKJvolsG8xgwrX7BBHyX+RMVCj4ep05EjyEgmzVIrI9v9
5+BnoysPxJHqCem9mX8gYVhnwFx4MmMDOgN0SYI4LcgMQZigtsJuYcLW3eyccCr5jQoG4cgA7TWV
mnyLDD37YaCa8Z1WnWwTol4Q8Byb81PibCp1sxvorgWmWuBj9NMlzJLO2wPQ4f/A1rvANetkqBuU
F1gOXXMXTfrmkaWMendDUN+R5enQeFS3VrsdlSORPJH1eZzOfr6eiLGhqrQ3rnHqBenOp4t0M3+0
ArcGs1qvkaivo9uOAWRtdAtVQ9sGL/9OZgNey/YC0r3YGTEQZP9fIG2KwKg3tELvmZFRCNeidnSv
R0JVcUSkw6NAXqAbY9URUfTMfbF64KOms2Chw399ZAr8Bckgquo72xrejUsS9DAdywD5zjEIID89
hYJB4VQgcWpPIw0eo3yBC+L5MsmH4VGkwF1yJJ28NAxB92Wkm07af4RDEXJ/dJNZhc23nhieA+0Q
katXbtvCdRpoKzPyMCzFpGkKeQR87bjU7tYKPM7C4TO+G6WxbVQXmw2rDFhWazo9kz9aY9hG1ROE
BKBDNmcPHX5u85Bwi6DWWX6C2iUZ4BFkXlEE5N8o8IeE2zGDUcAGW8aRiOSxrNoppsUMx0Uw0W2Z
XhcYh0E03ACd4p3SlzpXyLz7SVRWzwJX7s2G2+pDX7yf6CePsQ8RUoZMvs725s5PzbcCFkQ3mTJx
DjfOsyMY86kYohYnYn0ZG0UjGqXd/l7awZOSOYza1NmZKyqM5GBoTmokGglxMMANKCj6l12J++in
uW8IpHnCpbk1ZDy9bIEfDKbKdk5LKLVm9KqBV9vY+JZxdi5hdj+ReoJr/0RMcc4fXxG9KQ5QZCgs
jSbREewNAVEKkLe2Un0+639hr3OGT39opjCEDQvFSgZLiR4SWQ3X8+dR7ZUWkXyN53qaQHzfhdBA
ZLR/8Cr+WTas+BOCJsuv/yo3AoZoz1qE65owh+u8Hm+XDpAXBUajzuXEGyIknmzcy02XY3eAZUtG
ms0YsW8O8p2mi54jz+f5WeUetF65l+sv/ncMsezRm+0quleQxRz8GhgwpIsq799yfzHUPHZo2gJz
+MYgx0RUdHa9Os0rXLiSMd+knCCKcJaWpeNtfl/G/jGi960FOY+yfggy2a5xZfJJBts44Utb1blD
ti/qIKjREFFbwre2Fr3jTLMwi1xDAQ+orWV9mIF70wffT0uJyiQg4j4WlOX6du8MLt73v/2zA60P
W+efghQX+3OZGGYoKRG0V5z3ZRGCHKzxw8y7ifKfOIqsYv1B3GFJ6Fif9m5GWLMJNrGIBdZCeFQy
MVq5jfhpIsllCHNF8zksGsZsi/lKQTyhvFsbPlwHfLWc8bnmh64fZu7OhboopQ70gvsPrMOj4yVC
wEiDXgHjCh4/1ri1zGSqYFCxc3ir2YjhIaxorn4S+HZ1W0M7O5a5fhEakVUOM4UG4wycTSzB/nGd
vVyXSy6sgb1VFS26dgYBmuhFCY9lxPfPO9Gaq8mSIGjE4VervwQ5DNYWhSh4K0UnVHc0E1JzXOK/
vmtwsXefPDltzVFk1wvp2B5WnZa7Gc5ZskYEOtUcGKMaJGk+FhmC8S9vsTONdUqJDc8h+HyZP1SJ
zm2bJHxYI6hZJGyu6DYK9CXiUIgV2TsVsDFXU9i/x6ULztjV2Pkrp3aXHwL6Lsoq4l5UDIjilV++
GDzr5vixdt7PzpJHqBY+ZJcqkoAFNj5Q7h7Tjz6z0jPLiNGgsVaYHD3XHg0ejuKSVGzWNlXz13qh
cYhU52h05WxHWxW1YfdINpRv/rWimB9MhO9unSXG0kJftsDo4eO/uf4gIjriI619S5l2Q2qahnNg
TKcrHs/AYS1fWnthkutB5flGzaa2Djy+MfqHhqRtNtJrlMj9eZVRYmq5YJ+5BnhihPkoobUwdZ99
0CZjmHCXUd5QZXt5bhKqdPfnxUDH1/FWJ4MArewUurlFWstwOpIdO93RoqSYcm3R3tA7jLfG/Wi7
VTbnrunrgPBAJVb0ZgGgJM910h+8WL3Mjd68fb+mbwF9zsrntiXMu8YIRVH6Wla34EOTbgHWNDuB
koHCTttlVeH1M4vczjFa88xIKIS6Ctj1yIoJXorfaJejlSRtCSQbS+zno42JveGoCIDQTs+XtY1o
B15VvHgRPe+jgocskynWX++bnKh2crroLkFt1VO/zmIKpLtUr+MKG2DJ9GuzhfAhwyvihUhzEjyD
vuodt/l7kp5FatdO6++Hcoh65kk0LJBCvv2TWys/UMjymWc8T7HmXqJBZLhd3rSWbDG9IIEGGmP2
D4VawU2d1o/m8uszdD0tGtYNnHYZD1FS8hl4DYoKrAc7gC83Hp3bIqA3s7iXe2L4VOsvmAgKyQ+X
5LuTlqxGXEqMI/b/RvsADzio4YP1MJcsmaPF/fymNVHtgO7jioeAJU5hoMLAOgthA6QY5dxQBT1h
rWkw/VAudN2yk2u/a798biHPaN7uUAFRLJzhKSUsEWp3YqDKj8aXYlMBJLo6xpwJAs2YnSjkzqpr
E3xdFD+BSAXSBSR8G8ojQnCPKmaH1dLykkQA9mMzIvgRmLzgZnYRK19GmRLOP2BCcoGBtkIQbQQj
/wV0UWbyqdcTeBtq/1XZpZ4/VGLBjjual7lM4YLRtYfyaGlKklTUr/ECI1g7OhwJ8+0q9ejTKy6X
vzEEG2Ah8tyVplLKDYCVwd6aDtCPijqAl89WWzq1k4+xsVEzsndPjVVVemaiFlQlNtLjxEZen9RY
FS1kBvQ2sXAsO5pv1gSS9xdY5pWy/ePChCRImU9P1+R5IU6BvIO8Y6DrT2NA7q7rrHhdHhlkI/Aj
uwT4WNCksZ3sh3xxzLrOq0kYBQa2FRVhkx7Sij2nyCVISZrbiIHoe7LpBcCToseAMWAAyLwUDZ/w
4NYM9ZPJaQvO9Pjmr3qq9UJo+4UlKvq+boD5G/b+Bwe5RJfQqlG6HgVj9lSeHEePn/lt8m8muJ8U
dfoxgsshlBmNQE+rAWXsl+h2TbvwQvRxOPN+yy7sItH4ja+BwbyxKBHF367ULPefes6ViKnATcro
73D19G2eaVrY7Si1jtYAeg5O4qZusXlKPD7L0OOS+4RID4u3d5OZSNNWKA7bX71MPjGfCprpvf7C
94Sw2gMvBNCHYv6mbVv007nwb2RykAs5QmhZEVTvlUHZ4Q22b7hmnasaSoGiYwJwzNPHBGEeTd1U
SxN3dE+OgyvGgT9RhS1dTw/wbBV36YnkkZWpaHe6Gz9v6qkkZCRH3lVjfRdC7RAf62Jg4ZL/qpCf
ICw1IGEVyxfvY9c740ju3k0IHNa53brvcmM8OUuJPKknBiWcbjFlhYSUwmhuugns2FvvmSGPhZyP
eIl9y5eL0RcOBm3vyJG0/X6eb/aZlQ5D0lUbOOOmhcqLoSLIV8XaQvfgOBH4dutDWJMWj+8YLQNu
eIRXd6BrFGVXycTV351erHtypoUZ2b1xCIcjW+gaWseSD4iexuVYzFFRzA7/qWlMoXMIEfkHQTKS
sJvr8G+9ax/C5Tvb0Kcqz+hFrmvvXTH9XUHQO+XZMVSmkxkUymTnpbyEjcvHat6MIsmU4qoIWr3X
q2eCu3M4a1EFKIq3jGh9IqlZtR5gixkxBQdc1xsASsDXreGd+GeACia3HcTbYKcvs7mHpaQSuTsJ
DCIJIWZYwod4iS7icKQzGvdH/VqAb3caPFr9BbZCsStQOP1uCVW3s23zT7qa/wJd+ygOj7SEkeYW
zvlt6oKaWjMlkJPebvLYzOFJGmDt5OvRDtN2G3xjl2xqQh1jRThFPmXgzn8CLy8oyYZKeroqxyZ2
jxP+WamJoIYUm5v7AtFQAW5MpnWOMMTJbei7Qq3Z84rAIeViUOm2eT7OCtoYu3yobBq5H6e7ek1b
V5eOhTsTK1G4MzWSXRCTTHccqIiK0beXTXkRUnXH5AfdcL9x6kn6jgVaIJFMHOcwcxIzyu6znlqL
9nVdm5ZE2yUHf97OGsiVUiv1vmOJiwd+rCl3J4X9m2gbX+OCT02TK8DM7OpaYVyP8vPeMAcKi7y9
PyUlKdbo2BMrrzkKxVBZ4GktISoayR7COwNIyHZnIhrvF2BOGSSiDJwa7/IXHYTAYxSBq/8t6ApX
P0z68nSm1MLPWe0Yz/eD/0Iar1MhADtkhn/kCi6VR/kRbcoPJJ6bv5BPrwZiTCEW7jUsi5mUeFeq
rECKSejJFELySk9XVxIsU+gZdTcJBhoslQ3Rz3rY5KzcwqnS3YqoeSccldjY2eLZtdLVNVH9WpAg
LkvxuIiAFvbJaO1F/S/dY2OtLvL6cAf5GcjTPXagu60+kgIXazvw6mb8kDjZeTmsSsegzKfkAoMg
Vp3Hp3207COoEBPQqfmAdV2OpTbqVpIPBKs8q/NmQvlELrAqPl92f2OjKxZ2/NVhmfiPTfuU3Fg0
0XXKPG6yXgHYfzcJKh4iDj/0zyYriqLZ4o4wkUuXiTx2tZNCHgdZPBUhkyEgcTrZ9h3s34SzKI4h
jQ4q7FreTEBuIGucUHMZCNv9D29+1ckBwTAQe9d/XngdAtDG3jrTMFKCsJCotdiiUvs0ab6Zs3mL
7O4UiWz/wtcqKzzVItUFldtRubwRmE11yvcGt5wpQK4AiSkV7ofPGeMud1ReukK0v0vx85B4rqec
qc55E2xOSAv/J6I/JgG1bHVMs7n9sbJll9L5VObEJ7fWTwpci62uyHrP/FBtcfbAy2X71eoAHXsY
kAEMXkPPbYc7EPHCRmcROETkgNlESGdCT90Mpaqr/nkt1kU26+lM2oHVdqH5JH3lO80U2EHrsKO5
0Y+YO3TyerXHGtoO+W/WAvnMhI0lSg3On1Wd8+dKeZwUViIcmcRS3AbUy1SmzManc+FpFWBiR5bR
Ya/17jG78OK5jYmtju26/H/Qw6ss03326mL3FCd6pMlbP+5dbsqjzJZ2qTeA1p7NbsrAdlN21PN0
B9YIBMkaKbltIWIcFH6O5wBwoYTag9e9Mdgb6iyuu0rQ2fdTwmV0fG/27sho0rGcnv7rKAW3NLYv
nO3XhoYnKO1QIt/vdsnPl8NJMbcngTLlJEygWy07SP205SuxopPDTEXMOd4cST70gC1I8ziEWmVB
6qPJ3zEw/JTmOd/x5oD3hZFZAVqFb0BNWJU+2zR8qYJlYRnfH15c+3lkJ2FbtJFSJq2LhtzfJI40
PvotH9KUNCAnNe1l099shdNEXUwcXoZ6Z5xgMHuNBTJm+iJbYQpFdmFlOLgEabjDY1MkDS9oEcUC
1BobAv2Go3kH175VeFvm4PgwL7rj9r3UViowbaKJvOnzQ4XM/Hl83EEhBMYEkOHAQ2zD0x8ADQzt
swg/vwzcNY3MyB/Y1RAxfnp8uonQgTdc8XcOgEslzV5B9EMY7O4EwYCJ8iMJPL+lrVMVdt2hB6CC
WCXWU/fX33swV9ygwUNzF9IclkzOYArM+2iRUfU8DvqbnyfkptVyciATTXMNWlm/VQhsn3SEIepz
P3BfXWoj3JFW1UW9SNv8gQ+mo7poug0NaDRLsZMZmiJtREVGBddfcm9dTvdx65/KtQbncOYwBf4U
BV/Hq4lnCtTqdcXdi/ihv5D9WqXeHkT7Tem3j7DkK5UXr5dYCnIhpX+25YSKf4WQMCtL7edtU4bq
e1IHJb1Ym4lmJXPbUc3jxtO0WOZgo/z+QiW85g6mp3TdprrzI86xqCHgFM6s7X5DekbaCZZhvrDb
Xoq2NeLwzkIbE8WdIE2E151m0ZPgyhXhkXuhbSvajaFFJBokl+tiWsQ7RjpNXvBq+I9Ea+q+ENbe
WcPTAqzc6aJ0N9o1h27xKPB11hUgV5aTObOHWPll1urH1C0RVJbYZZh+uD1kPZAbXWIAwUr41dja
TVXmyDIODjmR9Onf+eZAlVHJEoQBYjAySqy6KgQasOcjc13zNs2bLLxq7RKGDapS3677tXTvuAas
DOMDTM9gCbRqxkWOMZP7HJRUMwy6VnmP+sMBPzXtiMFuNqz/kXlJwK2zS5rr58fMZLtzGlJNSEhh
taUcHn2h3wDG4/jO76rfLXau1PjZ8CUnm04ddyfC3XboRAUGiDHm5bw9gFLroJOCdlWxSkshXP7v
PID/g6UWhISkNQrywOmuHiEqZW+E3TTcYlvXsXYpziuNqDJE8Qb8LsKCjpR8rHJhItlLiDdQrYIl
YcrzRKEcFN2gxEHD33aLvJIHipFmQoBW4THEEBT00MIc999sL6J17n9cwMpUs0cw8JHe1p3jQPG2
FrS72Ph44nH47ec4dZGSuvvie3fPM3egPlq66jcppfHjC35U6UxMxtqmxErBCD6JyP8E3UutKa+t
lSVdidBmOOAQpo/XhS5pc9EEw4MS2WzyoxuWXHv68WtMPmrQefPKQPKHjlmNx7awv/MGXv0/e0O4
5QvvP+p2Q8vplwUUq/LKMaFDRl/4ODB2cWRanoHEzDPsh1X3EOAM5adFkDPPi2Vje6D+JuiKumA/
GJLfNEPmaklH1AhUvnpG9BdZ6Kco+H/gZWZR1D3ZhllWgwa2UtB3/w5uBJpJvCXQeRdr9B0h8R5Q
vUvLgJ/GbTUp60siCqPcLUC87v65aD6HyF33qjbqPrGTqrFSe9ck0u+sgP2bIqHTw5gQWgmnr2sb
NrSliFhN463/3hRU2mEALHeFl+mgQzrlt2lATKc/2Q5w8Nzdku9oI/Um1fAQ/o+5qq6h8Xbn+JdE
9M57wNj00XqOJtCwQzZ8BISEQPPqALmhtT4yDoF2dhWDZOinpWkkwlTZoG84TcOV2Lolgwwi/csT
rlT4UaBy3/Y966xn5GxXivgZpw6rxmzOEjkrr+3G6WE3pSmJhXWAUmtxhO3RUgIK5iR/1uHteG0q
qFMp5MvPYpPQAXdtQGx9zm6LUq+XkCQam1Nyal9P6RYWJbMMEbV3C9bAf/f+okdXsVha6Iq8eg5R
gJ7UTEFYBiebXbADfSq3fxtLuPfE6zhZAyN5bly9FNkihhJZB2E/In+v0EeORZHRWr3uT33F1KN+
Omfu5uo/Qyc24SFp/ZoFBPL8zeyGGpYV/CcBS+zJxvz/fr9q6ptqgY1JetlPIQ8RTL2jXzqR/YWt
IKk8FcANJM1GP4UtaBITb+yX9v7q6MLPjRh5TFVhtmXGlB0EXpge7o81n8POlkXVbKzjI43AwQl1
JL61GXWoXzNJLxgPc3f8pWTO1QvFff/4Uhn5jaDtdjODhATn1WZwHfUrWzC9hEGPhAEoIfwhFU42
na5yrZYNvj+khGVbtAqhXj8QbjjjwbLKxNFBq3BSq0GAcMxBilwAqxXHK6EKLEZODl0tKGw4mOTk
hITcXGXB0UBBncVd5vNO0GXUg9vGM7Tk1fwkdv5/lKHOMVsc9yGOXUjSPucPB8T0qY1i3PGVES08
GR98TTUNP21kKQxG3mD8ZCiSlHMOAPQVg2JDYw1XZvps+dFYwfHVGF3xtV0hTt+7VhdkfZUDs3bZ
5w0W4E5LAuQCvC+cCGjtqOXDTIAniFbjQ37CRc0J4h6LFuHUz4/RO7j8up5wy2S2hX1Awwla2WAE
hYNVM+Y3tkrb/9x96FV9ABOyX3VbZwC1oSEuJaMggtu9mkxGSfb1jxh+EvKDCJ+teW2ay8e7OfT9
8jeXlRcVIgSSS9co6mjF+yHlLHAMVNUO0GtkjiiDE4ygkI/opSTCMd0aKbV8qyAoIgFpTb/2ZSGI
omutj3CJyZ80zei9sg2ndrlHoFA5nn+CC+aTGt37661+ki0JDOisEPx3qZdzcXrgG0/djEoOvD8E
IsnnHzd00o1ZcRuv1i+KeuSB1Nuf7EQ3oVzxTJvT0gUGOvBhna9hcExImZAOVRgr+/03AmOUUJXb
rrDZn+6PlMuGcovMyf2AG1k64oa3IZd+Ucs/xXSusPAX+ZHxXflmV7F28E/FAPU3MUu+Q8GZknrE
2H/IwNLs08vyvFuH5V61hTPicz7QBtxYVFxAu3Q+z3eGtEeMZNnq502NkCXtqGwc8iLka/sT3RoU
LLIMTMZ2tNwgx+y2m52HmBBe6F+bsTtxBNlH7eLyqipI8O5ifawyHs1v8rMCdZPeQM1/pWC5SBHR
i3nqZQD0QJR2QXvOBQYoUiVudt82SAdmnBdAfVVF3TRoXzUnNSrdB4l3YMWMJa5hWffzVp6Nk6fy
YRD7NrZXliT5tnugSMoWfdkrRzIE9YrF8HozVICLAj56n/tmyhsT4/fiFVGfwZXlhmk2pDOS3jBf
wtWbn4QTEMggB1yPkZds3dc71QG8o6GYvQ/BerzUwhfpLJKiOD7D2e5OUU8MTwbvuWyEx5EJ9T2A
Kgsrq+M1TcCZsKQj87o9+reXdcipc+ugoZxdeky7QpD7dLA0QugEjAs+iLjbF5oIGv7/J4Wu+NUa
W2HhqR9BoOsub4UYkooTfW2u0Yjn631LJ3t2lusc4DEzQDqkjyzqgyGPSwxiUTx0ougY+wugCWub
ANFYQBHxW2kpBRCo/+TC0j8p1NA9elpiIXxRxca07FdTWRxYUFpTXYIWGcVYzUvepC7Tsig2G6dr
kegtLjF0tZSVl8iaWqC0SfP64vUc787NCpwDb6lS6dqUVOuoqTkFdWLIav18EKvKsqkoKywEA7if
x1mVvI8DK54Z6CoN9F23fQ6LkTqYiaS0GQ5GHQUKXodW2j4M//twXjVK8euGmxnSTX1hfXLEWPzW
eXsnk7WROh0PW+/6QKHg79Pe0oR2Nr+Ue5PImY23k4dqUmq3t1haJkC96B7MDEmoJoIm2pxZ9ScJ
u7rxQMD7+18dypmIIYLfXEt8PbpIMCubIZ21Lb4BwtocQpwoffs7yU/2L0uFqCv/p9LJh5DGhWhl
QM+vMDF8xloIaMJ7jSTEZFJKjcKUp4VKg5e7bh+DGf1NKUhaVkMzZj95yBm/O7YPsBtJZErFMTwE
aCzKhaQ4fDPAQUmN/4l6CyORnsUg3hNgyhyWJvZg02RJkZPz52FYQF/clNUOWOPLmX/DpQrPJu9Q
cpgBE9dHHW8sJqClrWImrcD789mGNO+095yS8KDdURFx2hvODRKG6hTRmQIrVyk4J76tHFvNFV2F
AoLrA/xM/fahokIyXzR4XkKiEB8zNR8tAC86Anr8EVrnxGspip26BHJ6KNJZhlh+7eGWDBFreq4t
aL8iUTmxGIxJ/g3OBmp3l2SCDZLTi1qv9BpbufYhbUV/K4zedsHR/5C+SZZXL0bYU4FfefyLcJbS
NYr4b8NNcQWoOh6v2pqrA0X5hq3e4axpf/g0g0rcwikd/rSMzlVvcWQvxPstr34VRicX8vDfefdF
ObvwWKDmMeS/li+XkAYqFjlLvO240YE5STwIKx1yiKrGqvDuKMmVosgKyKK0AXIRo/vQsjPUZe7a
lwARzZDUi84Wp51fN+sJ5SCKpEJS/wmKNDPUkr3my5+unSSlf2aHBARblO4ncab6F+3N46joasfQ
OSxq8dfFjRDnYMqpmdUgrxO5TfyQwdehawzRB/6ErKai9UwzAd5fDT5ySZJzrdUCblC5dYQU4311
wW12XHmlQWUnCD1oiwVjpGjJZAc7FFqUqEwHQFxp0aePPQwG1EYrCNbTVLBump0fnqW/0Qv/f8ey
Fi+nBDRWVBqR5aIE3o1TNoKqLNkwnoX8wX+xHWLJ1OJf2g6wkiuvK6NLMb62/fKPxotsJbrR9hYS
goAHgmMSEU92qLFw2AlrMcAFKAKpdV9g1CaLmPA/YEQj/B+rA7M1AozN0rGPrm7p5cGICWWRwxfS
mrqEk2XRZ3cjCWu71yWtmWtf8hGL30bBKX0b1/v/qyXlI1SxvfysjIFe+GoNCd3f3D4nrhqzbWon
YDCHtzUB2r7OMT0URHxqY7GDkdKzEt4iCjacRkH+Juv7EYvwo7RgaBJcWxBOP8s4UGJ5ot9St24D
U4JVHMtm1s1osMMAhF8p/ebk+ZqYfvizgBOd0yT9d5aFyuddBYXqMoRHRkNSPc+oX2APrTKcsBhE
H/djZO9BWS62of+MRBZztCTiHicOpQyKbDSPbiD0xH5H33uAjlVRbvPtSD8uqzQnA2EO2niGNifv
K00B4xtgvnROSZ6J1TdiXiX9drCyH0yZ1xAnIh6uCN4bIVzng3heW+HJElqbbjPEbPm4F7G3Lm6I
fzyq4SZxMnzrtsS6HEhFaALAPwXX59IsVrh+N0QHP42D2h+dwKowfuLJf1hVxvX91wk+tnnkAStu
M/EpnjUKKuCdUygV4JoPK3jB6fiOr2b/lNZlCH4UFESzwu1xr7RoKejbSRyCIcMk7sBmCQ6SYyJW
RS26XSBy6GrWvfRM7zOtunD20MVSuLd9Ftq1fyLNSzdY4UobnQyl8BV3YE2zjKjx/TbCCjbEMF5j
Wt/PE82FCPabTfcorC/AE8I5TPuOn6gHNnLTfLMcaw3lcBKf2X3y59/OrVAQIagR9c7QMPEm6W56
1UiF/ZG5KUaAsPcY/qiy82Bl9Y5lEI00fxgKgVUUsxkb7KhDKSEfSjk6OyJ+D/p+Q6SMFi30sZKL
RAyovhfvJ+lR9K3SeJ9ayWhcqPAzXMPk011wApPM8Ff36TW1+pvSBECokTlw6rAb3m99VnAbUEJF
1mShqGzvo4KuaWSp7SnuC711iQuGiuDEnKed8NmDnyrWnLug+bNK51yN4e/fVBsyBHD1Xqy1ovgx
pB+PqKs1AKiLs5M4vbU/tf6L0IZqd2gfASW6TrQ8OLbh/lYJ/UTrL8z7chdglXxbUWZQdJy67GGw
//iUcWDEiwtCCcb78Aornhn1xsaafW1BZf1q8SnOdAD6p7wf5Bl/dLEbQWqas1usYfcXLDCKVuUN
L0hFbXfNY6tikF/NoDEsNL9ISOVO/CCIqDCqNhyeIXkpayRvU1opsc2mt+KVk8Nk7qJjz3i+JdjK
7HdhukDc1Y2hJ1Llc6uljIbsw5DuOTBfEBswLW6nDzKcRhYNIHFJF10jHpFunx6lvj8jKeXHvQro
a4LP3Jav8Cr8gmiELeRrq9WmrVjjuE9ooJ07WnPIDQpaRccm5Ft9/I0G6KnRffvoYUqg8kLtV/8n
hYgzMa4+dSa3M8BKq243QFHA45VCq/x7XYu4DmyUfHBgQdcONamd2eqQA/Ws21dp5HoFvhT5/xNl
Ol4guTNKYE5KB8KO0P+FqtKyPgDe7OijVyhMXU9HwtkLhQimEsGSW6+LTvmIvkUw9TT3j9U55lh8
d62scUea/aoM2mTqBLmOpRc68qCp+6X//iPjyk43ckyg5/sGaHN5TDNr7M3lSYp7RiJLcL1xCGrd
T67ZGUZxQbw77+Ws2kvgvd/dMz8I23W9gSr93gRncbb36rZRM2f3c2uSGSBSJYtnc5IdB0UXyVAi
ksyNGUdBjQD30M0WEhqfp3ktDRNBzqCa4KufGTNlrThooOFYCwhsy+5t9PcVAE2WS5gsZPI9xp+S
N6AUG7vJa3S7ggXiV7V3UAL7lwLTYaB/Xh3MhMfYJEbLgarCR3UHuBIj2JODXusbL6mJvTECKcqW
d2RKKT3xOqfSiCl85c0XsH2zPcpzk+tpTBS1IdxdVTiYH84DHqjpqx5oUprlsB6DCICigX0xG4Ep
2YljKseLwAIAubAXFqvLW8g7Py3W133oQAfUVhUYLPfPtTl5Nda7nBUVCQotI8ukqIk6lNH6R0fE
aaDGyCcWWYGwv8EmK7fXNb/tIXPoCOX9xH+xLw6E635VZvz42f2aRATfszaDzfBuOGYV6PJfO8Gm
cK78knnKa09Ghl/d0ikSiVc57av23TEkBDVAl14VL3EDcJmej6e0RRfZhDl9f9CJ8GF4buQv9LL4
6r6vEBdHsze7YGcPdOVndj/9Vkp0SQF8HoHJankqpzlTiMDwSuPX2aQPTrlPF/V54AACSBlZv/59
b90+IhR0Y9O/g6rG4AKp3SSe5hn6zbNeWEK/0wF41J0dF2k/kbljHPT8U9B7jEBm52y/Ezw+ER/J
N1KnV5BjpJCdvvmNtVj65ksUxdb4Hqv5Fu/RPfABu1bKIE+bJx+Iod07GioAIdEd31HOP1dr8W5g
b7Lj5r1QBRtMXJ2CBMuaKtGTEo8mXcRSJ7GZU31DEOI+w7aZEF1SDbJFPC1Rn+XULWLhClmZQ7ZQ
0s8nWs28fY2Q3E+ze6cdZ/BJJDWr6Xt/Asii5RI5woyyPMF7D0eE4hh6KMOZdl3036i2nHr87LRP
wjgPd6L3NewFjwfijUAtmTL3hfjwm6ImCq8/DxSrbrN2f6M/KQr1ayiG9S460T1ho7V76eSd9t0R
I71qs+f55sIVfupjZRv4t+Nikrv60P9GcAQxb256o2ZfdcSbeFmobo0l8mhdvzZH3DFA6fds/1R7
XNNtiFGFUuHDK3T13tSp8qJOfOmuVjZMGvK+kHAUnVmIkv1ZU1vLHlabZEPsbOMj3diAWo77a8Om
XEpsaBRj26dxZzeIYozwM56kg4ZZ8l4yCwww08pTE+5jvKZDVmmkroSz+7Z5XuLg2RDYwmV6uNRt
3FhOMZsxwL3QLrlQihE5pv9xew8IhZj0N1QkVnoU6DcAyiyjnQhNApW52IlX7GZYzmWPC1xic7hZ
/cRhtxKhRGkyEkfyJk+N6OKnp+3vy4XqHSbAjqlim2LnPgxQ1zDFG+9msDXG39eZOpi94nDtlPnK
LFMZW+igerQmdqdDrhKtFdrHRC5IhSou/p6ZuWxnAOvy9uv3MHp5jTziEiMVUUbk5V8bmUOxwb4x
/U53Pu2ZZA+bCLBviSQMbVPVK/82/QKBtLsgdhq+lQoLB5xq6dO3sMKMIpfchqSogHZQ77TJh46v
HHEh8N92x9t207X1FfMMvjz3oJPUingb/zW/xjJJKz84539V7Ktu8t68LofPWSkBDPEvqGDBqXxr
zxYbY/VnIipfGs1Bh4EDkqeU/k/q3lXp/qAHZHevnry9Fe/aOdIpkk7ESWwALSaXOflDzNojce0T
7DfMkgey1TdtLONru5BOO+FC76OLJLZuS209WZqOJ/T7IAJYpnsaUuO7ltYNOntemNAaEy1EbxKi
uSubZksH5B8cwd2uZrKpawr5OrAUmxneSinh5T4XRfEUkNE2YBRxxGFOj3mSUWyou5LggjPro1Kq
kY7AtBK0zLhTkQxk/xSH/cr3jjKbQaFLNUbTI3bObABjpMVSKfcziwm0pcMqeItY18lwqNwLRscq
zfn9rbhrv5rsLMf+fhd8pRVDWSombbYJK08yifrnYBFvKEHYIz1TLkYs2QP4TRY1WiCCh/7UJVXJ
erC5L4MpLHxQzp6788Ishf/qWH/0xkOBtgFp8zJWuEpFIpa+KXkGYyyqVVthaZvhIbcs67WhnhAG
6RINDj5OOSvSeMWzFKgVTbQ+6T5BipLR5tURHqOVAD7G2KsVuDqNhrrNolY29RA0w+kcersApCVn
+SXQE0Smhc8RVHbdSdEYu8uEyKYuUJn3n731svH7t+wgI8DPc/wKbUd6+hD8Bo4I8kw3WCxO+9gO
uY8z1DRL0YRMeN4w9/P2VGntmnt238aBYScMpHS6VDUd9I/ocwcxWSCodQ9DgKgwyQGqYILxpkiC
EoeReQtZ4cznoFu3mrXUzuhQhJQef+YPzfN0qmKgziaUE33HQCG0j4SKnMOAF2IjDiSJFcyn2fdk
yE+mTGi8kNiY3doZCAC9xYtFt35jsNCPcQk0U6B9zlmJJ2gxRbaDSoPdKD2/TV1FTGwuiE1neJkv
Gjer2x4/rT1nOAfus2aoXWCgPEmpU6JHMIW8PUgyT9ks2KHoHys9gUuy8e3+bZrt68rOhhGbcW1y
daodhyX8hFvF2MSlUDyIUAloh8eDSolhsp0OGW1ECeHRDsIvfZbf2gVnRc18O27jg5VWRL2KhTaY
aut2MpoP8v1v10T1j55KbbetFte40nEqmixve9C/s2zdCk2cnVaMKEFXmpUxHx4j69YoCv5KEqbC
NW7KhNqFRbH3bTQvmbxq85UfY2rKXt+Td3l5sEq2pT3lwfOvC5udwDirwmM++CNNnV9T91ZSgsB7
p1bucGusXVZOdPqMS3bRuwIdNCduuP0cXDTo0hxR351OWWruMPY84dzcMGKgT0j8/MexWM9slwe0
cjEe9FYTJOUCkUWhGbZ4G6K6w+ZVzv/teGSlqVA3GEjDpWGiHddvx+WwRbcWFouMKUoe5fuVba37
S/nMFkFl9PofNdrd7J9lSBOsaU25vzeKI/nShXm5iSNItQANYK0gOCk7Xi5osUcE9FkUFIHAILID
GL5w37bPynBmgtgRe0X1ajGLvUuJXvJGmMES5gDrQsa+qhHCYc8HHtth+XFBjeDnRyt4EasSnION
L1dMgUPV2hlhetEvkoEAdh4lBE37lDNLgfZCURpWVIVz4LgRkmawTV8/YpDZJjRxqwq1k0Vk6kgq
pNGm2m9feLtr9nBKBazXe+ITWKMyIrQJ1oZVKRXuSkTqL+ykakGtzi08lhMZU+p6ysXr5HV01Ld6
mU7hIKwsNc3r0f/4O3jXgGdFDvNf8AsxaDjQPb7YWGFSUoPtxQU/kI27N2WVat47xixhiWx/R7dE
lb14RaO3haR9L+Tz3jWqdTJ3EQLkwXDIbOIItcU+VSp+KaEpl9F7PD9/TC53qIV8+j5aHgbBKi5p
bK5414CQS4t8BF6reVErWlVUAaRVlA6pZLtPzoG8gX1Vz+kC98zZOHb9EmMlotb1T7LJrDWZwcc3
kQdYOg2KTne19WJEsFGnaCjdH0GCX8fj5H4xoWSb4uGFxJ/l0wT6uWTnlqyPI8iXcT6C4qCjsJe3
F/wX528PIDEshnzDm0lQ4OkBnFRaeQvkQXip4wzo0JnDmmKGr+IztdFTN1JbgKpEsaX5HttPSqmU
+vf18+ZgFhsbvUn/d72ehPl6EeDRduJO3XsCj0blW98MR2zXupaZ510D6qPwRokgbPjU4VX6QyNw
5S3hFyScH5+r7wyKI3pwQL1odVYP/eI3HBc3VhntVaJwuBP8rYRDm+JXo4ftc2BPspl3yJEFjUIF
+zOBLlQKNT3hs24MeRXe0SRuWTP4ndUV+L4ZCR0ChPW5a8mmm0dAK9McQONpfG1EXXlgedqOHIxd
uc8wXCt+/qX6zYGKYwAYvAreP/bNnK+R4SDvQSL7AiH7HK9yH/Z3rDDqSlEV3GWUpYXqaozidLMi
5D4Sb8RZb+ot6eFRLHJOx9JVH366NCtl9A8OrP/z9pDvUqUUbNgkupQ7ymeuHpDfYEeM0bv9nPSV
Nn/PCOSd+ivIyUSSizaqx+NWv5Uk43FS3lWOOQKz7Ju7K43+vHy0ltwbQcum8I30npnz8le6a/HB
n6LPbismovPeITV1BVc3iQFPTV2eqoW2kawmTrN2yv39/Joc/SkMnO6vV+nWwPDSM1VC9C/W2nFA
AfXZdcS4SAqBdipx4DM666DSyNl/t1z5w4f7dN940ZZ5U+OoFQ3J4eNti3k+zIyaw1uaMX9HEtKs
4VCG86fUn9vyxPC8H0bebRl/La1mH6S2dkeHGfzWmo+gDA7Qjjhs4RWy1N9Uw4g01pNKHhZ3lOAm
wROlmviHYna18Q8wmOC9oSkAJcnceoxINgf3jXdqpKaq7muQAjE1Ol8vB0kdU8irF/KVGfU1TnwK
b+twvd5dqrJD95OgnZ4mXD/zzMY6XaH27K88cNErxQ1w/pJofbBmH17Zr2rHdVcrQa6odSt6zST9
ilKim/s4eB12rOeSM09yL1JX0u3Juoo5vnyHyi0L0u8q6/fpFesnGqnacrEXl9N39yZmhWC4AAYu
vTHu1QuPsSQxtmrtbxBBbStdXzczkSXWN1rLbp/a4MrpN2S7U4VqcCio6say/HG6El56MzbW21zv
xl9h57XeZpMIZxh90fXbr9k/jlSWHX5yt2ttyenRb2Pk+BGiANRRQLqaphu1iTA0ce7IMYgGAXhS
Db9d2/zCeu/BWw54JQ+o1/YC/LZOfR5ZMEbLcNGibkEOfQmrikmtupJGV7X7KjHreLWEegNrQxJz
ATyQ7vKr94F59hnWTDwon8Bfx+pC4NW2igHbZkLaW8qprari7WJfi0VE9oIWUGbb0sag+EQqDLH0
nDQAUzzQ2XTdxEbjQnbgrAgSt3zsL6FzUMfBo/ZPxjAOIdxHklwsQz4Yn0we5mG1UPvN60IfxIXy
tJnlq1QmvwDFfbfmLO/OR7ZOm5B65DtgkgpimO2SH3FFhElfRaPf/CJAbXNOKXwTQ8vU/Un4i9m4
vT3thhEOVA4w4DDaRt36vGzPTqx+XpAVoyK4d/HFqEUBrLpU52rmUV4R/UCb2mGC5AOnydGeCWgk
4WtlWjZOE2v8tWnjlBfVkWkgTRRb4XZ0Csgi69prJ5LCkR3DljE/Dn+a4QK9U7sssVyCuE9FnuY/
TVi5GYcrYm1AjqKFtFcgjQOyOGj5PBRb5QhRJZOfIbqD8ehoWNDZhQ/tIuRR9vAtTRHhePxa+GHJ
glfnNBdGD9ICJXWFrFPfOOXWMJ916zKOeIrlVf+dMvtiMLZgMMLP/NRLbDPWJEGZfbXp8PUrCy+b
/s+cJn007SbckhOUQUH4NOGJN3KCQkgFGyEmEynkpv1poE0hRC1oCVug70pGuYg64KS17lrtQiZM
AKPg1MHoyS7rTG0z/uP32YmTj0d7P6htJN7x4/jOVxSjmVT+mFFYPHt7OYWF0cB7ezabWnkb00iB
Zu/3tjHAOEaEZv2NI42yvydnLkH9kXGN1zbC93V6KZa3N8fKQa2G3/24PuSIWIy4pcBIsT74pnt0
+8248Eelfzlv/oxl/cNUm0fpyvHgjsgcHMejEpupVoOxw0XM1Ed54kyFJninlX0kkhH2gXbJgrde
W7ZtOfLMbPH3D928ukxxNdD4CY9MWXqFNAbfAQ691kQUj3P/mZyoK3wXb3bWBcw+4Lhgug9FbTKI
DF7Ns9Jpx7f/hT7TFFe0jX4lQwMjQbaSzX7szA1DqiKXcogQ+7pWecR+P0rV/BJHsDfvoKTm8cEz
cuMWYBomrMbR2+be2J1JzZv2m9hoBbPEKFbsMphW16QYNLN29+kKW8yB05OktKGkz0s7/VAuAjSh
7bOdVFhAwsZpY82lPW79u3iZ6ibWydrjJYD/3pifQo8h+QINpfFam9il0Qbel0KKjAitLGvxJkFP
BZ/KThjDeTABB8JC0UABvNMnkAXysa88NsdZ6hBgBD6cuThd5UcRBTfdSp3hzaiopfEg6+KcoREV
B9E75HhjCgQ3dR7cjSEnrRfCEFCd8zqaD+ZB9IZFGFz/Lwvu9VgypQn1izl/fQ2jVd5NSApyWfOw
SU88TkpcChLVUuRMf8FNj7JKAYiGDwLBWPUbOLzq+0yXBKtVVHu0oeH6ZT8lbBcrBl4Xp4n34HEE
SkuZr/mWdOZy1Du0GJhggF72K3cqAMakWTwkY5Pj9syGUtMK8H0Km7mX6jUUWX2BIPODFhX1KGvV
bAHPcDuhTJ8NYMpq+dPlBumn4fayADmKGlSloPZbboGJ4KpCZ9Gebcs9CYEOMMTo4ZZFuVhZkHQb
tOWDuyWXNhIKwHlHcyqw0BPzK8ONA205JkBFf5lCNVHvUxexKPL6Z6ju5j2ywswbkXfd4j1x9gCM
WP0syMGnP1Kh1eCvKOcm2f6GXdXGtB1rdrfW1lukNTvhndhUh+9EeM+2JtUa1xOjOzqMsysmvlZC
9I6vDjqlYKa9FOvQ2BnRb/xUV3fQYSR1goOU0Dh2NAQU0qme/tcY4Xw2q6dlE1P+ZYJyiBOPN25+
K12+rxk1Nc1+TUztY/beX6S6HAI243qUK0mpA8ZkULF71gQEONhdnUqsqBBd/iqSWJUo6bGQ41iP
nFDd7Ae3wjz13ByTUI89bU+EATcfxSSzr4NFZc/d81meAa7DhC2kt5XG1JT5B5M9OPOuPAnzz6KZ
Ulwd19oSwfE7akxCx9XQ+BCU34iGhdTTbbS3RUNlNGupKIGVwEFSsaqdAfJyIMCg4rtkBnQrTmBe
HTzqDv5wqc2awgHoDsB19UZl79dc/lnF0MLUVjc5ZhLr/2KL1imjtlSdTyYCOB4BmohnNMnBxXlJ
I73TfWLKXJsOzQD78/iKDcU4FKzLDRHUjtCcPFYyCDnu3OjtL0teIy6AyuODhvsjGooZMWoidMyS
qFhp2Z9jv/4UeLHtJxswDKVua7zDwhR4AJ6LRqfiC+LJcotJWqhELR1Eu7L+Jy6pJG0YB3ncjUI5
qK3vRERmrxfOkqdPmKq/ZgrUaChikhMNlE/a+Li4RyvhBq83dATmNElMKMUj3TDF9w9Wn5ZRTDaH
Vz2qm0j6Sg4bFp4plE3K1BDb0uR9xZxfK1l6PM6tiR6AhPlSIVvhVqvqKgmdNJjdVB0astMSAQK4
GrREsoCK7VnyfKVhzak2xteakXB4OCK7OFZRorhEJr2GY5xrDh4OHZ67s+4SAnFmsgER1BCuWwu+
xI3nawnK/kyxIDSi5nJqRx2G7dG/CpbiGe6D9szIdeuZE21ipVxmhnbQUvmQ+cph/OKbAM9aY4FP
WZT3FU86Ei2OnsoQHPuKc31iGxvN1tvqzy1RNSfr0oweog+Xq0N1iS6yDQN9m6b6WJjvimqWEoEY
rDn+uSeFN4YPccqrmfFTaHzfX98QBIxOgrTg+ASXyGUYS0KMZ9C7UkfBbvPkRvayqlM/D1O+XL9S
sNGMuedpp9qeyGN7180x+Q4qlIAx2H7VKE1ucczDLlOShC3qp4L98Y9AOT+2W3LzJqhpYkU3+m13
orU5UpbCDt/5SGIXpCi0IWyFjSegMEwkBGOfH1CJzIYVb3umM4OKVZhDZGJGcylnyXa0XXbuFDw6
JuREbj4RzuzkvtvXkIpJZ16tI0hKDBOm0W/HOIKqIc8VQqTOA2eVB+qnblqzc0why37MS7SeaFk/
GoeLx7VdzMTvzbFZDJc1ZAkgXlgHrGHHadiQff1OZOlM80/Pye+bOAvcBvyavm8T9CIrOg9h8Hr2
RimgZ+xPi86bo9KHxkfMXIUq7NBV5G0kauxRg+x1Q767s0AH8MXUUFdD0o1+aB84sk7JQrjIbmnd
2/du7hDVPAS37zmPz4mgzYCg7l1mtnaChWFH6ZaTbEYtR/wuNFab0eQ/pTS/Y1bf9zLlbBzBmtc2
QCsnb2Z78epFflZkS4kj2Lwg1T5eTNqfGbb9OgcIUtswdruAHgjZUc30YZXW2fbo927trzTQ7STp
OGeAwQWj9wslQU8jsLb5nVv5GMZCC39GEWH6HPV+Jj+6wkQVeR4/0U48A13VwiJf4LKB7h0rxC7M
DRFRCjCEOXyHHxb+1QrSaje+bIrja3OGlCZCXpjZaZgPNVH1Oqbo0Ag7z2XWzKM0L+oXRrh7BQ9i
WhorYMpOQRWke5vchNnm8J8lakMYo9Zg6lo9apwHpBgOmpse643nkuibEDzgdqcZyDTQXYXBjk7q
4O/Y20vh+hIAEeZ7lQwtWwIbBb4Bx6ZR1I5SeNCSLYKN4JHFnIpjaDgzOlXd2RIHgEl62AezEqiG
1iNRAujIGxuRkVo4UUFXxLFjNfW5G7/0hsWUiLo+KbmpMrKp0CPJg8HKQ8orEp4cBRzT1Q6MoPTL
Uy+SCrAbMqIjCk1nlcXR5FkpvTpPyAjYA67B6peATzXu+Pd8C5MHIUZwpGtck4WQ12hrAtePBQnO
ouzHxQZUOM1HkVAfjX3PDBw4DbMg5WaigvonMxIzUuVCecp3FNbRFv3NP4tSmfYNncyPwiQ4FJki
H/ID/BgmErymJmo9mi/VClgyxRlvkoemPFx8hVk+U+vC7EF6KPgHFgqk5IKxFpRwgKQSUjgPNqmq
WcJLQmRLX5RCwY6jbLmQfN5o+3k2chJYSvZgQQhrw7q5Ytg85Yl3B7DIEosNndtYwy41p9MEuspJ
DOwBAa0nzSFmjrr5aD5NRZN111mkMongv3b0hdGEWH9/N4c2Eqv6wSJyVp/pA4CrskS5KnlpEER5
3D3M+4tTTtGbU+oRZTlLqNaKe8Y/Srr5/rPAihFv23q76373snSukWUmJ/+SeJ2Oxgiq/gBpGOEj
2TgoObzjV5Zn46a14XUkRZ35ms9TJPYjfOon3mU9y/LfjUfiRPaGhJaLdork4Qw989Z5eTuiRT6s
P6HDZT1CAbD/kOVWfpqTDh+Aea95TuWTPwVf90YsP06uWMPBMzB/yJVe4iX5TPI90n9c/1epBcuX
hMYv7ATmPRE0ZgnCBxFAyBPmqiZC7fcWl6Dt+bafhPG3MDhojz2vzoXy0PWYXongR1ykjJoAE0e8
eyaY3vpk1aMkbzV4H+ItrPfk/TgCdWwkOhZOVMoVfPEu42ZI4EltLil2c644nfXgJU9aQXmUM+vQ
hORxLyzgosnMkyNu2oDlMBqycKaAArKvebimb3fd+rG9VxnyQQckhSlrwnpvO5i8a24rO/k6tJbO
iEQTWyhNYJcEBqwc38fjWNVhizk9ZmWWUvX8+WLRt01B80v5z3HsWh+4UU5NLgyqnWKZgHRMZExe
Ek11Pwpo9QmpFquOVniNYFobCWyKViSAthIEZhFPWafW+/yqqhWItnX5LRUIG/xP17mV/EsvtPTB
6YWuIk99L8zhPvF5vCm7MAcRBOFnDeKAnojjmpZ/7f0RKwYWP+IGaRxm9PVawA93vDFSjTZ/FYHv
QhV2kgOfvuz5zMuGDk+skGQW2SVbgeqmziwsJahKHkClLpClEg014dWQlgLFfmjSwHqQ02NxE+ti
CyIMvA2uxMfbDRnpoNCOZ0WclZ+vcCr4drOlgqnSYcx3ijHNduC/HnvIaQJf7AL/GkOt3LlCa6tf
skL1abv/iG04syeuHHOkApPsfq+yGcdQiNvdMalJ8Elr8tI5hl/gYEhKBjzrJ4sGbiyXGpGt6/+1
9vai182V1pv0Enna2y1V7oi8xUY5tgfx+iEu2QbzLTGCNhBHbjqXJEppMZCJt/8Ah3xC7s5vunTo
Nj6sz94TKD6kzky3c7KFUSEJ6QtaEMpQ6bjXeRP50EPDFlK+KXMYSXNHH8THx76mB27Ow7XVPuzA
s0wOL0itiPM79XbIubrotrzOTRGBUXNAQ+Y6P932ne+RLXyhhTGdcmHsofHPt99+mp39dbQoUQ9+
8sql+XPDS2xUhT4Jcv+rbLRYC0biFhKvWW8vGxhlegyMuyhUE1Vf8dTULUMO8OWePYG6mPrOdbAU
TEktzqv4bQ6IneJDIq5dN88j0c9wOOCwthNAf10cBe02807frnlH2Jz+oaPvuihPEakvfwIFbCj3
gfqgWT1TF2KDquUlYpKndQth3xUpIoj1/JyZrZr4rmVc+f3VI3FkZ0duxU+i4yRy+rqUh6qoAIyp
1yESl53u/PpFAVFykKoPcKrp2BIqoL/FVU8QYNFS8yggZyJwPJjtlNAmsc0LEyqM3MrnMTxkm4VH
pV078gADoqfkLxcWVrH+U4OUM0dCe8wiAHbdl+oxmScZeT5nC0s7Ix1wVyQLsKMBYedl9+EOlBZk
WQHoHfFp6DyhCBW85xQalFpekdt2ll+XSUtOYm10kLGsEbMAJ+7VMwXBIl++BDngjkPQgeJkheoT
8Mao/01Bobvi5/fbzJ0fzk+ZyfwWaQxVBpZyK/J3zLM+q5m5vtcyLzWpAh3/aauN7LcEQ8W1ngQh
Kpd7ouhhVKIt7SvHYVNJdqLpGHmdEQBodnPjfN6O4CvvXwFd4YDQMfZ2w85f5odUMmDXQAJMZ0ur
Uu6JTvXCl/iBkMCWesjSCy2i5hKGi46/OifABja3fbMIZSJ7W+xiLZ20uNnZ19ckLxVHH8meqGT8
uAL8ZTtyQq3VVGqXRVM7ZONr4URPcovf+e6Z7buDP8UUq9i4RfeMBbexX6fiY/b6RfZ+8N8V1u5R
ud77avr0SurEH0lvk11AoFOX351ZpALlJVlH0MzYOws0HnYKuGyzB3TslrcpjrOh//aDoxu+nZF+
ZOIqEBko9igAVSpr88Kvshrw56Yh1Ihxb9I7ScazWtnWFC3FtoyPxtEZPe5taLEl/c7z3DsAY9ft
BDWg71DKTJ//yNIsvhmcjKsveH5PkhnZKOjIiTeyZtgqx4zVAFJ1egbuf2DxKovdjKHxTq53T66w
9TJn9qB1fUlNxeC3uM2vVMkgjWfqkvJQemF1gsp+ObNNlxrav4Fngci/AqaDYS/yA7YKvugFPnvB
TaljzOM2dHkqaqbgn5HlHJ2viWIZTYxnW8iUI2xE9lpokt27AHidZTmhVHfNb63ufh7txefdsfME
CQowRbKXwPJ5S81F3RA/ScIa7z2p9eAp1asAYw9t3f4c1pn806DKeRmWUgXwc/lwI25PrETqVeGT
JpCHdl/Dh1iG1n/itpUpcPMApMFZF9er1RnCMqDuuZ624BvuxGmeJd/NM88/5tfgNMoFwPe1gw47
HkJ3NRGx4yMT/ZifC/hS+6iT45vpaQxQVIKAH+kjasDKqJ6pfV1YHjY3LeCQ+JrYe+BqWSNEEBjT
csbQzKNeiQwr+jS95iseFTPVMrxG2m4Xq7zlOT6M8PXUxLrKbPbb3FvuOnsrD5ywAInP7ctC4noW
AqYf6/ib7ZQLnwTubNweCkNx1ytyqnWkgEtZMOM1jiMZ55/flStqNhkfxyJdDcyHS4VptW2vEvji
0XWuFK4VDJUWqB38+gfAPmOMFTrPHq8evw+fVDJzO3X7u7cRXwYRRzg3yFpphTVSwHQmVq0YhlWQ
qcDBgSsnoJwdesIhiz35uXfyZGm2sgnUmDf9ykHDwz2UuinUSlkzQkFJHv3II/554gVKOuhFTyMC
TsmRug+3OGXzhAhIY6wzHq/LNHKghFPqoPa1Y6gLd8I20TIPwpMHU1BUtIk/UXxDHQAKqUshxOM5
hHNR/vT7D0lxQ0TEO4NT7pI4CqqF4F4JvTvNNca8IneHp8ylG7fsGCS9JXH8uRxjXNvuuYUPmNg0
C9/zvgn0WE2ck0OhWDVos0FafJmHs45peFwSfFFSIBtkJd2jjb6BH2scU4LkpfHLOSThq+T9iX2v
mNlrKl+IdcEOtlXBSyZYRxQEo3CON7KsrF+HpRcs754li0Trp83WGCbKfXvluUNwbboARCFOLvic
YRkYkhYVgMCW60tQFuZRvli0t/xIlwZwUb1q9h8kYsOIp20GoV7UNhB3SLgn1aHYXgrSpLeTm4Sj
gOORqrKArLQBVbLBDfJB7hNuyOYADC5BXcJse//oepg5LvFjZ/+ppPjj9JR5rYN0tjUDvrZuy3xP
YOxD+CEHGG50RzHd9I7/lsg/TP9lgbO+AwuqHzQ61sbh1FM8yDwMUg9tpcu/VV8ANl4cmVrMpJLq
nnlFp5RRc0L7bAD3GiyNtVqV4FYBJfN4DjfA+s+MZ1lAqMbus4DdQ/aalXJN2SMq2zX9lQkDVVNH
doe+oM2WnfrCs3lBq7q3aQEDpAk3nl/cXDlsY5NX7wOI128xKMuNfcaRG/Rv5viQOFgiL3MmCiyD
gxDr05Ds8HvpG96DxBa9dbFvgAWwqRnCMxJYTkew6H6wd9ZvSXSIGEHXF7OR5672SfYAvCB2a+Mb
sNVx1TFdjW3o3qfdPlLOp8G216KJqBRk7X/tgaDSVWVJkvbR1juAk47xDWBz34nzS+m3N2Ovj3cp
S+00pUigZRjrd9qsys/J5r15WcahB2Dsx/BWhCMzCFnfV0IM9oxr9soefEkzYL1FKdvoknaAQTxW
SqHnGGfUnazPlXl8XhIkWS/TZb4tkdl3/ghrYCtJAY3a0AWQSzkMFoFOHN8ZamY04lL0Fz9BDxtG
1GwXutvCzzdZktVQis0vOH8JM8X1zOLtZ2wSUuwx/Wls09LB1vs68VIb0QwRU75wfMftagZR+Eo2
lRb6/W9xqx3NxzKhXn5//vMZuPujM0HsiwSmPZMdewSIkE8GuN5liEl0zvuPbXCAKsnbB6cK2Vjd
LWhUgPCWeY/Tr+HkZrvwB32BQ6AYO4OYa3+yLJ8IF8CjiA0Hds00RRFJF5zI6WQFsiMPzNstI/Lb
9xqrSgnLBcHMUluotKz9WIyvQp8XD2ga1bmFEkvdg7ZiAa+RGdLUKuBxtJ+jBDUW5hwLpMZJUgiS
PMNulNRGclihBNGOTXqdcjONgDRLNStK114JEnUuJd3WjZnpbZc/Hh78y4WSMJ4GaRLDvgyC3BQG
rtsGm9je/9SSX1ty/+eJm3xQ84s+l+3s78AZjBq1Y/2lR1kQV3nN2FhC0trILCgtucXV+V1XEH84
ce0V90HCzWhOwM55dzZVH2soCBKLJbDmQbB1lMnqTATc5nIKz4CsUdN3Fz/u0O9NS4W7s/GbY11+
mkwKSrruh46uXTqANehl8QAl1/sMy/zwg349os+48LchCw3MHRPQY5p2k6YY10pohWXTJm87aS2C
IJXpyYeUvMnVKJWUN51kM+aDQbXPt2UMExZd95lsqHgxbn20uAcu/uR9NmEjpzBOhoy7NsR8M19L
a5v1BCHbWehD7W0YT/DC+bNDfhohoJ0teesJv7w1Gwx3VZYNTtisIVQ5sCvpDOkSCw1ze+w4uzeE
8F5bpahXyOLCf6LAe1ckQOCavljuvzNAS19af+qAE9ZXvfkEykZJMjoW7T1p4vgcJbiTPiDndJnu
Ztz4WB5znH/yFl+Ly+r2IVA4Qw3WNxZvEcBb6VnfwhpjAaJFkonjy0oAtoZrzIaCEDPZ93pvqqw/
fYLucI4gFdigmv0lQUbXI7P1lJNVSfNUGC9QfZxKWG7IpFVagGviT5GStZ2TLZSIZ/GeUxDo2JZJ
7XN4NTKltsvuyk/SYFFx3U69hgNxNBNlfOxHp+csVJYE9CQVy5pqDIueaRFxaAaRJNIaCWwWFGaV
JFbR73tPSNb9kbJgkCWPIWYAIYw7h5QecI9JNg2qte+4+IgbTKRjT94KDaa5H02W+VAx6FgDZgZW
SuGmbMbjibIFihV/Y0e7+X2RNYg63i+4xfbRFULcJDbcR5GAzPvahvUbEsU0U07nwf+UNGCcM2GZ
Jl7ZwuIUZ9r10n/y2NkO++G+qAhbZHCWBYmkgx7wnNPyYz61CrxTnQLdrzmlwM8l7HCHc2q5sfJy
N/TeDmFhJk1BvcCrmD5Ff+ktXPUh5WHe9ve4h1NWlTYkN6gqLnC+IMeB9nXGXh07XdRKuq9DAH6l
YR7PDWnj5W/WdPTodB0muEcelEkOf8IK+XaeNUZgqRQp+QWxN5hhMRNBApK2YYeKBgETH+gfuX0t
34w7uZnhn2oyHephUsMtjm6UAoeuIU40iKnXbmvGyrRrakBdgBPo1e3/jXjK1kMcVTa/E+XeYxYj
1oWiUTWDrT80oSCjG1bITf5aXJRF/rpx10gcJg7j+N0IGEKWDzka2EQnqYPUksuM848LIWiyX5lA
lWgbSoPdMkK/ocDSsP/HPtMFeSBtTmU0qV0Fl08/gDTCW3FwX92zo6QLZVRvIMCw030hecYJXk3I
G4mIDt8CsYtSQjP8w3W190ZpoZV2YS0aJL2tnXBTRy/xek+yoDHSeS56nAPO8/pDc2VWtllPh8km
MFMsgSBbOKTr4UTVpIAxcTUR/rXHmms/K/BRsU+umOhRl2FwoTtiYhuF9n2KAlTOEwz5zDVAAfPx
/tQqRFKx4hI5xa+RmtcTCOHPWzysL6Opxj/V34wqQywWg84c/2ZZeZwGxGNiPVtPF0Vn3pzMmVic
qtNEF/7NRxNK/BJSR5yZUJ1m3McYuQcvMtMdEybplwJIn3CMmfPDSD6a5u0jTx0ADT3Z1O1SfbVl
KSKW9/e/YW54IKuSrk7PihoD2JLMDi8m/kv0v//V83AX+8ViEZBew1zq2WI67fcCYoKEa/EBzppl
udGRuYfaHFD1YNrOsuotgp53rk/Wn8KULFJUCMsQnqNbrQic2f5M6LQSqehSwf74deA1Mh5V/ADJ
Fv03DEBlK6syuhzNN++sb5hoSYbBS7jjBzqnfFLdiT3dOUcpHIKHC1dRACRhUZCHuZGnLNn82Up8
RoO34oEZpR1iENoBi5+eoFSnSSP+4JQrnVucG+gHBY5DegraIHdi0kCsRf+yuP1KBa2EtLs0zZha
rHaM38VsV+ehp6iNooXUwr8pBODJI1lVpLn7/z6xf0Vq/zbzz/+VhgQLMcFou/Vm//5lo2QnB3Pi
UBMIv2qYFxHweIw2tB3F54TSrNgvHt6HaSzt+itmWS45mvgVjcmtX3a+w4eUmF2la03BYk7cKXHD
ukOAhYeToxEiDvmysjke/nKoK9ePwiOyU7wbPn915QkEbR44FNtKKHk1lRiv6e3cDRYaasUd1vJW
Gwdyv8QUEmOozwl4YL1+jNj5d7/ybo4HB63RGa6Jx+sbw8Rk95BsixcXgQpyHhs58XfyC7dfcEOD
ptjUk+xVPzytXgFG+hTgToUuNuobj31sEh69WZOZ8KN6HgriYzQrrSqCovXRI1dMO2OnqLofHium
RmOSCM0w8lkqjwuk3o4Ww6iiixeNvUqYiq989rztAb7ZTlmvBpgd+jh5nKTVKkSrIvNRGczLMOSi
n4JWJ3IwZC7t59DzLqKgV5QFzJoljohNexRMvL1z6OBTjfAW30AYVGVxU+p2koRntT0aCTzSizqn
L+hxNkAxpAN09SGaM9JKw+8bGOGP29DzyguQnyMcXewOPl/Xt6h3DJQuR6cxyU6QaJOyXYSaKUpt
fRZrllz6Yyq0UvL8oXghfrqnGYLN8JXy14FEIp5XZxe/QXkBHlnb99JN5aUI90k20UIgBpGJbqXL
iDVFsoE8b5Ir6GP3FKLiMUEccFEfvmvVXdTYIhmHm1qY/O8GphwHw1bVB4gfaNW0wuEgAKgMJDI4
Lto6rX5cjmIMNCh2uJCuT7IHMcPFTN3oiDdwaPA8j0md7jLOQaZhKD83kKiLqMGE2qZe5FE3IbjI
6Xxe7X4P/CnjPi8nSCankikbmEF10ZsUCYDx8eG2b1q15wFhHj+FLPYKjiJA2fofj+VFWTk7EEFv
5NdhSdH7BnMfmr+TGzX3FeSGV1tPm67Xabxf0LGf7MuTXh3sS/ghpUwHNQzxIs/s5ftIZtPiZLx4
lpyb18vi6iJ6U818mO+y4XX+HA0lajY5LEwPYQzfpEjOGZmbexDG65unuKzlPn/5LTOsZGw7u+6D
J75/jKQ2vjy8bt5pWHFMY6a4LE3mB9OVXE9n8FzmTuY8yol67ZbyhqYH5B9UslPOsmk7EDQEDHpw
2rx/XRksM47ks0ADm0a3Aprh1STYbctZ/iR7NIbr2M3HdmVbOoCLztCnLzLHP/LYdbR/nwfuTtLT
P9cpGDK265/5Ak9QA9yE1eBrlpOwbceMwK1UtSbKwTbgUp5G6wKHDOjvKs9a+IoQct3jXCUZ2ICX
uL9VZ70f/cBlNLbr18suZvqqbImBPFJIfUBdBM6mlKL/VIrzqJlt9dDZHMNrFQSXYl/Xp6o/Nmty
6sbG/j1zldISwLSs6Wx4Qrqi2qP6thiiLDsT/xk/bojuvVqtXBSF2oEycEnaeLKZmRiQjuF/wyKk
VTwSbCnVEGCgptCcpoez6He3q80cUrx80EUUbSS4RRO7hGLS9V0o/V2MMkiGCgwfeNgNsBlLdgwv
fXbbG7L7UDkSW3rUnnyvN8S/HazJ19X1kcgeWfMWFhdtQxM9lFIPdLxtiG2tiInoShr7RIw0o6tU
twMR5kAJ9jsqB9Mlrilrpi56t7aL1nJCsj1IGVYGxyIos6rELroLjRdXCvSGRGrON0LFJ3gKozw/
ax+ToltBF22zDs63yzR/0XtWFkAq34ZejoAl4tGy4jw+S86XeYS3DvWekE0DZdjNQxtO6vdMR1rM
RJht8pzDqXiipoMataNUp8QDmQp9iXE/ubmyFGXyZ6zoSUfsjosRlJgpjC7E6lJ/dFzOVU766AVU
ydIdpqI2vMG4UwBTdUJfhzrjRiW2Adn6BhxSjnMT+W221WdEbpjOnHccnZsn6lx8LvZEO02jN/6E
zLLSvUSfxwjAc5zGKEf1MJ8DxEbaGPrKXRncpIzmsDRGxN1iLOF4BONCEvm7Q70wH+25BSE4I2wA
hJrcQRi6Y4o0q1WrsuSYOLGKxp0GCsP0M3WqCpP3P1Gt7RYl2iJiRHQTF0u4Z58Xkt3EkAbzLeVZ
tR5kBxddQ1ws+LA7TKCEm1udmK/lhzQjA94YTXJAugovv9ZGYLcI7+8s8Z394RfbmwzzMv4O0JhY
j0XSlg41VL6KY1TFxvE207PHUGyTS+PZBQyTnqA7CHMQlSqx6HhdpSgY/wMInz5+8/KTxQW6u78+
yR6sK7IVDaOiIOcL35n4NGe9I44rwHFAEotxjbhiiTelxpahdf2ZDKoXJ85eSkknbGC7BTEKEbW+
iJ3tq0PhPjGZ7WhQlAU4+1KBpK9j/3TDiWusS+EBUDmdcEhjJUI4T7iO8Wv/3bAz3trvY40NJHTL
gHLOVkLmfYGFT8dB0+zEE9YXu8g6yw7ITvIu76E8V3RwsW572M6Tjnx43T4a94+XRAwtHsg2gPpw
ZeX13/RQXQk2VsuVG8pWqxe6KE33IcHkNeUM+W5VHfFRbEqyUFuW7DjADuCUBfI6EhiJQsWqQoWE
T6V5PhKeKLkoYwm/OBp6XID5R3y7FiNe8wANROa/2VmxEjMAXfIkmGGYtX1IXWXb2upbkeEsHv7r
zsX8hEs1TK9nC9iFW+eBpYd84W3Z15UpKJVLPzNNuQl2zUWsvYyuhhwQp/vHbdHM1zIB5ShcNqbT
H2TyP/iK/L4O5xYX/T1UUhWmMFXy6FMgB3D+aHd7t/Hq95o5c2BBQdv/NznNhAGpusbVJaEm0qnY
LTZpvP0q0TPLNlpqV7dSGD547ztR/uyGOWcTg8RxZVqx13fLwN/afKRuUyrlckPzkgCyc9N2MPXq
CFnQOVvPtZ/ehJKH40xAuTR/LAnPnU/+6pHVl9fANsdAhyQLLLESADKtV+NB2U79faLhEw5qo0+l
ck/WKXlGELZXkJXUdTtIFs1yb9FvGeEcziuURZ0Ev8QD0H1FMFj4cFnvXZyxnhXA3EYGYiew+udy
btCeLwOaOxLBC9n0EVahM5Rn3LcUBeSs3GPQwmgUuTZFMkAxmXduS1l152SoD3tfbCv9/Pc8hQZp
jHQnfQODp4uT3EEe1Vime6d9FXpW95reK+xPF8u9zZH2LwmS2006BJyUBgx1TXxtiKqII/7xDX09
X6N9eKI2zd0KRfBk5gFyCVZ1GVzSDJCkFQd+71cuYBIBGOookr8sBCWenUHnJBj3cjfsaZoAAc1b
grNigj27fYLseFjRB2GOyZDdCrBs+ZVux+0CRDvraaaxtFee+dff+RbQJjggIKtHbxsfIBhMs8nH
aMJs8y9v2BrYfmOIUBXW67AMl72hCdgoFRsWNcqHZw5ncU3Avrnm9k4Z3eEfC70d9scy2c5cFFTD
+W3U8qqXHFXz3/IlWgS8dS6SiDR7e8XQ/DgwuMAGcqkYVTKFYmPB4ZGpe970129EOU0l3qJgCwp9
WWURnN+CVGBhoC/805LDVszmT4bqCBrxivf1+BG6soF09/C64OmQlnkoc3iDRqdmd19QGvwXJ69j
RX+xWl/DASpbiuTWggq1m/duq7XomAvKXxpCGmvjSn9CYf5t3yHqihMgqkPkSBRhcQrdkoQBI3Fe
6L+WxE/luYQGO/BlVoAevFDwMu1pidEgWof+vUHOvQsp0h5MlK54A7EBlFYhNyyEQL0RwIAO+USh
WKy3lB1fzo3D4cMOFJpZWSdlwHLZobMuc3oQTj4Q4kb9lnzyYnfFKZd+dWAHQlprPzmLX52nPPI+
YAWXk9fSgAi2lZPlmCrTZZkWqscyrdTqjhjByWfIVh5cKxNQkByRLI3OqA1l4IAfOmgkfVHsQlZL
YcEDX7yjAX7GgSI/8STL99e2LEBIYKnqd/PG0Q9QJWSpbOvw4KNNBbRlA9+ldE8gsJw7cNQpTCVH
RzG7WDeE+HKVc5mYtHoRmpjATv4FPVWpUAEdGHiN9Xvg5abWfdJpEOTZYwDENaA91hgTQozRbR82
+Ndvhy9ftuyQC/7Z/n+gWUbAhWu032ogwOiDYflnlZdjR12JlhUNNSYcer2tOS7D76+ROZd3S2yv
TFfhie4n0YYPFAI5QjMo3VdQ0Ew6McggM5RQl65VC7Vfk3vE1n9sQTdfo5gL2ozgVmjTjaqQ2TfX
iD5lF1dP+pdnh/VTxJOnvz5FFpZJJXcd0o3VE2d0+lZAwgtM4miOmkJhfHRQ+ojrR+rSOyr6dfLf
TGD2wELEft4RhDruI/b13SqYDtFb7VqF2ZjK0i2tXE4eAQLDya+zAUxdQCyYCnuv/cH3lGzVaxrs
3rf0plzhc/EEAG1Y64KNObvR5OI32YAaVROaFEyGMZJEMIhXcCfHdogn8tU6Ci4RG5g9V8jaO2lf
Ncb59I2Ve9V4F1AP6uxR+OyhXquoHQnKaAiCFuzB+B+Bl0rr1LDbkNT3HPTKVBRGKTaWCoCy8bYy
2VwYH2q6FNfrKyUkNvvJp7rLocMy10vTC9Q0ow7Us2Qj1NTrST8fqJG5ST0NXdb65rNvfJqVzBNu
MGYhpVrUWIKi/Z0jhHavvkpLJucdYQQzb8B+T/NJolJ96KQ1nKU9FGsQe5dJ+pPVLIsUWbUiQC7q
JviJBI2fAhDJeWZQSBxyU8gaTfNl+dO8gjeT8CJmc5niy8ORIuSkDoIIN3wp2qtYBWnbxPzQZsse
jWNWh0Ka2ZxCWqsHwDd7+5SxAwv60jB4VHZcCFh3b5tjSgHsysbNj6bEl26hJqVA3UM4LfIVUl7F
wNKngZclePg4mSYxguEcctokMcgiSu/ZEBMctweYlNlhWrHADXssEzuGuxxtQ4gWvkhWRuVanSI1
D9An8Jn8v5xHrqqFIL3Zh6TadrVoZ81zw97j17v4Hk8xlgSZqNa2LDj8gXc12BEyWqHjqlknoBbc
tQ0fluWDTbmUqgmGPvpaAKsTZUVHNrFttUaZeCtOyW3GidctI2nQGpDngRFrQ7RCAu4g2/Ll4e0/
dnhc+MyjFUChgwDnSVDGq+8tGoi0J+RpBRJwVcBX72ebWZpVQGooCCSmh40K7c4+mrojyfWmV71C
q/9O/zyWlRv+SSOfmivOi/OODrMlMNW76aad+1OfHsN47bewLWoHjyq83ZQDLqwuU/cYZ2UGVjTv
F1Qv5zIOiWlqBrzJymwlSquoQSmvRDhVSiCluZs0smaxxMqOKF+XuIRPb0DXUhtYFvdemxNKXCBn
aCJfWePrhTwiH+pw8yeCMnsbkZA99gHd/lKij03M0D4RoMDLffdUlwjT/WdMzo/JGGWNE4v+6uYl
TnGgFj0y5y3fvPrn3mkrTGJDKCCZgN6DmqGAXdbQBsoHRhqnPpiblbOAQxifDjunJizriSDUbr6Z
43AmoY0X6N3Y2ep6Igrpgl9ZKQr3VCKs93bm1ZpO41Hw0ASgjO8JgP/to5wXoHQM76lC7jn3rPIv
M1e6GQ1DTu/Vur0YmT5ljxeVe5XfudPkkvsWKXDLiDwXfky/XlumFOYivp2HkQwjMehmpSayM1pO
OXGkL/6pyg4koajGvqGNnHBjVVIsN9hg2NK1n9BCi+lARhqHs6U3TVG2azeQ82Gz2nbplML/h4Ub
CynQMVls+EiI360JZR6Rv3AQHPOJ3acweAzm/BIXUd/UfCtkzCaY8EmFDr+Xr9b4w+2/xnEPg9iK
ivvgzyofPXYfA86cP61tLZvL9xqg5JDBqyXHTddItLWaxPcg+tNSNQ2rSw4ED8i2RMgk3nJ0BHx5
bFlckHOb32m00m5VaTzz6rGLyWhSp+Oi/p+J0GKe3+4BbxOazZ0tD91eP2kmZuU2e/hNHoqXQ7JR
fz5/qi4qmYDqtR4tvlxhf/E/NyEXKGIIvpT2GCgJjqAEnvjkOvfoC3zASijfHVnauxDip3DDSngV
EBCMlOnlG9J6iho8Q+K+A/2VAmId4FkB21MuD4lXZi907abnadYQCSFgKYX8pQLX6D00dARYPdwk
YaW7ZrtjEROlKOXIZJCiMgInpKhEKcZczzu8b7DTp2fyEjX5t0Ia3lr9PheJhlwNtjCrsABZyYIP
XkHvlvKUxY6FUINyqzRBXgyXDJbAxMR3FpdqfJIIM/RVxXkfGp1xqRzkW4QMusp7z9kBnwyf8G6E
zQGlItW1N53drMpxr0X/Vdd0h3daaWTzclCfghTj0BNDq7MTWBn1uxL6PLIC0lkVZfGAtqx6t4y+
rE2iH9fBXllqaI+dQAOF0F6kCKDkvBRmD06Ettux7fjtG1NErJe9292IToAvDvhfd71Yo3JWcjtg
F5QC7Zf2jPNceCppJWcjLxkybYQo1tjLjU0Ckp+NrU8UK2rqKYg/hRby3maw/YmJ9Ha1G7UlxB7X
Lt0JwqW66nHtf0YsplCgbSHwcu7jW+HNEpHmO+ekN72IINYS2vMzQBS/gd2NUFKY7MK/eoNNgkmm
YECvjyPz2J2WI4nY3l7jAc+HjXjWh1i5fQ8X16S/sUo8V6HjyicEy4VpcavT/qsNAf2+p0Grj59Y
ZiXMTlvYnmeerlfrWND0WBrwRHh6bHsVnV3QVmcs2nEs8WAOfSSOIjZ2eH/wxbYctl86b8EStPid
Bck8jxYepaR1gArhNrN4Kpu4QzaEkRbykCfTRdWagRekiVOkQEr7PmaEITGsrG2Z3tTyaJ92d4RT
FIbi4y0NBknF0iJr4loFuyH4UyobCWUMnlIDTF0/SVk1X8oRuJ4fAAYUA3Kaby8t5vHAyb4AlTnN
n63WODliweOogg/rwiLwuQmKf72yRV+84+1grvVtQjW6EtnN7Zw2HJIGJCXeFz74Ls4FVB8z3+JM
SlCLYLbEBvA6OQG4jVMkyrpJAOep8V8QgQDlBMdhfe5SLucPgi4gnm++n5sKhy2eWWNq8VyXlASu
+xngrT4FXmqywo4EjPX3lw2CcDc90B+KWsxJ8DAv07fgVJzXmu3GxU++yXkRevSDdYINyWI6ABQF
u8aHZ8dsf9QRRCO1BaUEZftD9SXa9d0P0WGjlwCPYsUH3VuZ4Ug1+YHGrjKsPHhYIC2Sc+eOj05v
Ze5sXtXk///tQs2iDsneJmk+SbuaKWpjeaWP/ge6o07Pnt3dSwstpG8zR0c8LEz1Ebug8Ff1H49r
7aUyd+CAUF7/i/KpJP6Gk2SxacNVRTt75aCVxTpme3a+jQlLS+tQ5I8u733RvlTYkXARi8kdmk42
XEYETlydGjvOazUolbqFJ+fbzKqmn1RsvaWE/TLXT+SWLjLqCRJBkLM8jJgPewtQzYuT7NTn0/3A
XiGWrobvktaDc5LcNXDvfjMxuAT9YX3Iqx+HaILPGqAZ0KkLOCSyUWzeCnDdOdCSjJ795VV2k6C3
vwEhMxW1d+Eq6J5xm5cos6zvtFXRJht/zJWScrl+kHMnWj0f7jspssh+xSQlhnDgmv+5DJvJKCnJ
qknKhiKO3btG51o/HWfXGbT817F7dkdM/CUMWpHLdTZO/xGaDlgq6V5RXiQ5A3e+qVEy3hq09OBg
4lGFi5vDKYfQ0XJGLBYfbqTEiV7sPcS2faH5rGB1qN8U0I+JeQvXOXhZzcIqpnCp0oFk/Rch/Apd
BjiioVGaAgPodL+a/wDD6a4jyxb9oJld86XQJEnjlstZC15xcw1MEw08vjPs/mNyOamZWH4lveFK
m7s72kKJBBaZMomeGIogzYX7SrvwyH5GbQQTxnawtr76NDyoSeoorgttBmKZRqt/uQcTdIdqPFzD
79+kw4IceOIDACqrDgtaKrx/8t3KuZnyc/aFs/FDM/elPmWaiWLFHIbmWqFQz3oZLufLbo6eNxPF
qvkMXm1cgLfFZJ2bb8n+y+2uftVk68Yk0o3d2v/ojaMvETM7Pt09aTenp9wD0kIo6fJRZ/XyUa/Y
QtD4/q14tlntAnk1YxqrJtn4MbyB/eJfLcBhG1GyqRF+r7YfXERqdPQliXvt5v5RCsbkUXh/Hq0E
ks2+3tjoYpeMFeu+V//cylDlCmIC8jDcQPvjh9+4NqYJ2lu02hV2WmpN3QyquqWAa1uDfHSuhAmo
gAl5b70v5sKRcZ2uXIiAR3hvUCrXYgiT0aGHfY2k6nr74f5VCyAA82OM8/B+yDFLUF46qPlyebBK
r0mA/KJSvn70rYnXaEFe9gZbYVs47J3BmRB7tHtsKWzTTkBoyTLhP4wNB5iQ6FB7YyiSt8W2umPu
U3QO6jOxbTCU2vECapIdWyRWHzu1doGWBLnQTkho754YuwoSR9NG2iXrS6UaNdVZyBeWAn7KDJ5M
x7xFv0gpe+UFCGi+O3sAhWfw77MN26yf69Cxk7suWDD744mKv4YvoPhs/ZIUP3W1bu/72cMyZeCP
CDfZW1hZT6U4muEXtPnK4QNQnEsxqUJMtBsN8hGnxbGZn3kLg/KG/SHywaPbEKsXCHSSfLZs9fo7
0qt8HL2rG/JQu36FU9BPTZNVbstFLh9EaN2izyZ4Fs0zLy/bR1OM02Yn/Z1OXTf+Fw6iG4NdrdEB
RqjxeMaSD4rcptM5kgxFm54unwkBqOTRv0SLuyCp917LxJBluCXsbdr92fykxM+6Nyw7VbX2zvmJ
Xyia2vsX5i4EWJ+Usd+7SVq/IXWefCHopT7jn0DZmrdGVkuABC2pQn19vvI7OngIXdHFP4c1LVYF
OTFv9jx7g4M/GcXZr7WmIdBGytXJFMTRInnz88uHu+5nTwHxzq/gws5b4+AfoaGS5PwsGL83M3MP
fs6Oyp7aXtzW07WOJJptwBpd7mIvc+035j9jE8+k+Zh6d6BCo5Bk3hW/fZTjZQeKGBg+RCzK5EeH
ECw8NA1OqK79Y2+zn8mTZbCubi9NsU+S2utl5/JzTbWK6OErJFue4gTL5E9bmu17jYUuGGIvh6tL
HUPsWdfID1fNizF2/fFztB+umrkvUnVZPVle7atVr1ZuKCW/Nd4aSOjbpeW+OWgvRQj53WUad93C
Djkg7Gm7iycxzD97oAynNxv6iUZ7dML8p/Cn1DQTTIo0LM0a2d6pKOUTzDwQIlgDicBGSrsfb7NR
KFMJVuli2RlK6Q+zt+5MQudPklXSSk1KpexcW6KXyeGnMK0Mb4i6pf8eXuyPt50UQGUmCvQ1fipS
iAGQVJ4nlwzH3SjD1q8Fk/gvI64u0M9SAI6OVTWLpCXD+2uoh4k/xmX3zKsB+b+r5vtdXYR/xAyy
UfQKvDZe3B9RsczKJ6Zwlo1r+foHlYjbG/jJ+1IMX4gbJDFqVW/YMux07CYvqEYLITG4ol0CWrai
PjlyxYPp3603TBaF51MqKCImRIRtVa17i9Czb5J3UudvYgQOaR2t+3nOoa2Is5QyWEfQxOy2GQg8
15apNgIELXse0c37gUxl9a0D+ETPj+9EZ0CwVKuZktSBktu9y+iqYTyJa+047HzbxnGo1dXJbLk5
3+os6awQ6PFYISDMPJVHIe83nsVg026VrFKLuGTByNNJvVETewkXEM9PfwrZYqVVCCXhd99jdDvg
MtZvxw1Wycbo0ryIu5auKqk6sC8EWI+TYfdeV+5dPxyO64QAMXx4Bj9Rl+r0jnKyyEfhzLGrVokb
GRztdgnwwzHUFL39Ubo62nWj7dhDHjsK/NF1Us5WA6TQ25dLy7So7v9n60FoR6RW84KCy6PHjiSo
T3gwexc5TkFKN6APz0ae5Jd1mhfHoYbBKWmzNplbSoybDsPjZVdG6g2nGxqvdzQPWGvaokiCbDJC
6EADAaIclxajJhKboNffGtW3ROuQdR1grABZcaYBWaY5EHWhoK7h5H3yZorsjluoaaYpjWM8+0NM
XNX0NTgSxvWILGwppR8vpTlqn3sCuHzLzQ/fA+GbA6+ehj1hzJaVADOi/6omEPP3Vyodwddu7Ooa
DRuPfSIfilz8k1obM6m5WD8j+3yKgynbj0kq6Ybp7x/Txg3Oym4xIsfwrJg9IKuQRrJO7jRu+s11
FkGnUNv1FvRLNFxh10+gFi9wE4XhZ267AqHyLB+QqtqCCugZJnfnf8Oqhz3P1q6PEXpzXxYA7kS4
c+zKJpodbhu6iu/awrH5kIKyNHfrDcC+kOjZ1gCAEkM9a64IQuuLp5PQbV4r2P/yJBy/u7Vp3kAK
+zLde4wSbqDCoELzujjdE76AWJCg+T2kS9t1SsQi59Go2cFveaIcPJWrXLOUdtSv2SPBE3T2oom6
5ahRIn/S93rrTEPVO1mq0xP/ZPB/vX1kcX5nzJYamyF0JqVzbtWqtfX/HoR2pOGNOxDgaUZZbWba
fBiNHVR8XvGQBVvfCZG0cTrrMBInjNpVO4mRTirMfn93/B6aZ0FFqtpWcbITn89PD5C3T9iodvM9
iuXAhNOsTOlULG16Pa4pyODBq3kbFnmNWastJw6WBzYjdO5AdSPJaLVQtku9s5GGFnVobzXuXVGa
ClJoYk15s08yS0yt4cxsjce+WHyK9LNKNCiqy5fZVSzQET0G71OQwPCqEGbIs2PJvTGlRpraXEJC
PnLZ7b77i8yx/YHrvoj7MxLPyx0PVmR0gRDPkuJNKUqIzC3qQGSV6IjWuSQmHQQELnxCG5Vy6aoL
NIfe+0bCg0X+YVubfmK2VguM3YG3BlQ5M/DjVKs/vBJozHo+zTI1c17fXcVNBFZvLZiPXLonzN4J
525K+67WoXveA9s8EN27gIhtzgG8cbRB2CNr3P9sWQfy0N2zlbbtqaByNS1juQB+F4XdKjnw5hmw
T3DSUnUdsaBAklT6IfIWiDCyGyfqQRF1kYZDdBFJjuHU1Teozw6j/iRlMMvlBSUkHlERVUnUmlBZ
rVWafGkDrQHQifbMV0Mu0U2Fnq4FZkUrU93rvgCZzY/E4DGAlK+8IaTS2wEa7+ZGhssjzTkBmssP
8yS48hGUUYUObDDlwJiq+8dW6pbcho7qQ9XYekfnz3WbCMOisimy9Hzhy5lWPNTQn1R1JumhTMTj
U9S/qh7R325ZKJhQRxYY4lsXiICifpTztOHKfhv3zZKTZ9jBOx0eS99Ykzuu8hDwYQI553crBt06
WK7WeVFMnDuNxEsaTjZQMtygWF7p2P1KzUUSm0B2xD+K4oYtWjfnt5uKpewCImf09JsGmrqOJ0zY
ikxOCUfS/EeuOd+Q80qw80ZTnAOiVQ4WfI9c0/f6puuue/KLq1Ct+RYq4O4CFJBEUlCLik7jDGDf
eehvRB3ra2qEq7WuA0QsvVKobelVlZZgDOM/SmcBnJs2eO4/hmuVBIP8s82RgbSC+29NGSBfGDs8
pimNyuAlkFunmylLSwLqK0+e4ufLHJENzmGI96JCip5vhAUiqU0DwSqktFp2N/aLkk19kuyGSTg6
cI+eF014K2psAT7YdxFGl9l35+PIkgOT2rZuAxhxuOw+LV1c0Gtjpx/J21RyKqbhaZRXix9ZMqsZ
UDmGZYzXkOy2wBQA1iZFhQAYhNu2UWA8RHyjB65FIapQyeUmc9aFXM42d6cWd/z/rSzh3zAgrVRT
hjjBrPttuLXYAzWgvTvyz9qRepaHscRAjZQikbjuLs7NwA2T/jJS3t/qDngnwobEiADVImIYqP3P
2TQkYFWCzhF4DlC18O/qj3KFmHR5fhT8CZVA6yWTT0T+PLxnpizDK4qPLMA5aPsT39D35dol0hj/
fHSq3fGOMrgRUZKv5BCJS6nUmDlH7RdCe6ColrNcBtykHF8gbkc/uegK+NrUycxDQA37va74QXsF
ZYnDiJyRfvgDrhwHyaBwKmRvMBGCGjhljepyq33GdbGqYQ6aWm2h0nvTUH9Qrm21djCPqXlzfDE7
3qgxjsAF1aNUn+ye8vTdxG0uqWLXM3MrAvZAYl3IOTEUull/3xD4rexaQTysOv6x4pmdgLdUVBBL
DW6/CcHzGr1cFrdeEVY9ybZkml2Ev/ItfQQ2V4EXesfyFrcXzzAZF4Ee5z14E02VtuKM/42xbfYu
51r61m3wruCB2LF4OlzsLLGD7ie3dRrL5Hv77sRwTVQHutnhKoBUd31m6Oyg/Y8qYbNkmWbxJZvr
8TUsy7va0OyFfv42+LhR6BpC92C0a4eO8g3RyuA+fcJuz09UpaZVljH03vV9Kl/aZWi9Tcy6UXEB
4EyARI3uWJZWKb18dAR1S37g5oQcDd8JBeP2XyKOyOMD7auGfSYMcWgIj4e24edL+IJ5y3E8gKXt
5HjiQMjq9mEa/A+e5rdtwg8NfYujsDBw7PSn+zE3WQz+B/wX1V2wIOIQ7EZMWHZ7g2zGXU+0s2Pi
CpVVGoB7VHZcDZQHFXWkGutyFkMl6lIKNlCI8jJIgqkOFIpw4cv4Nc55Is64gmb99jwVJF+Jc0lS
gtNVUI3oJlTH4yfbgsSvrwfZ2JeNgbS3lTkNOHd9xH/dKPXVY0T4Vm4DImdoO36r/n5WChsOIPrZ
+RuemPe8Q0n5ixlWsMLf5Gq3rv/KOdAnRYVPwep2jJ1f32g/JiDr6/ZNWqKkB5AsVdzqIhUKQuCW
VUOfHvjTLvJmyPJkEDVPZG98aaO1B12SvbqkRtQPyWCMt/thHn06GXSXvdeoKAhmbvpVQ/bZUf4D
4QWP4A67lJ0JhGBGmMHoYNGSaDYio3NEykZSbiIXN9PcL6SRHUoi0BIVCBaBjr5gqLU4HJefHbfL
zKVFexiiSdG2zzJqIaSm+DbngM8ZSF0SPT4SEkPUwzjiA2PaB/8Ae+Py2V6aOzVTktog9pPo3kpK
r35safH77T8KLOlGWjZxGK6zETz3dIp5vhhx91+qq/rGQEj8IQOSq3t6YFQfCYDU/XeTQdcclDam
NV8GD866MMk8H3EFv3xZD9nVWjZF0xyPgTpOGCGLxTAQiNyDXfeTKg8klcMYeT4tfQyCZUMYxrNU
D9EYKeyQXp7OtEbrYxezgC+FU+SePJrnkOWN2irbrhxDw0gn19OM9U5pE9bKtIkEymsGfkejI15V
aGkc6yN+34vd63S0KHZAF+ocDBM2vm95sKdmSeKziRWHpw0HVfOHfvfhmlesrQC3NsPrB2LSkhPb
ksB8EmNiNNn4kBcqXial32Cr+Yj9x1lhRLMfIfy+Jc/7Y4i4bfwXMJHvMTBGesEv6S3ibzbVJ9qB
CAosLDFQs69sHlaVphNZE3Fjw12WSbxDZ13dM1kgUdTAfO0YyBaMuGsZHtct9Z7+82aJxzAB3e2Q
fg8wNbAPHJfKBdKKIdcHW6PYWjlaK/fYtJnIo0FqpbR4lSNlDaaj+IEdysiG9XPnK/mKT4iRioO3
bUrPBmIQ/brHDe4sMVBk1WHliZZRzRPOaNoCHRGS7DpHB4DmkVmA7VsIklEVbyYf2X9HNlbcEN5C
S3ZHnB6nxvkqK+ZC3WzQ/bYGqxlTKXjjaUcj1BNQfdvVerTYAABXPUuMyRVUatWLaRDidUIW3uI+
VKWM9jneX/LtzvX01izspNE6zni5GIyZjTVPMrYuI3lounXqBgDjqUee+48CNWOR1mUawxJnOSr1
6L/9QlKoM5MHvFleHuYVTACj0U//UkLjgNpJLS9/pA85L/aSz3cNk+LJz23i2whVP02WPsnGbzaV
QpcVIEkybP85L+R3kgsarma6got50dyTQgxjK56lZM4tdXuIHyV46kxNsaboWr9lWQajDYSGNRo6
eZSh/lIfZEqH7xvNsTkwkHC1kDvAgqZ7cK3rrNJ0b1rRdsKlzZPK9MZdFGxPPH2pyIzPS+KJaxcu
HMbo1QSYAwCkD0qfUkp6IB9spDFon9D7K71g7gd7jGF8mxi5W/Kn+TmUVPbFxrOUKpepzHvKSxLB
VhFYUrfsFBGaN0EjB7sM2ptkB6R0AIhWyQ4CMWeTxra15AouOOdDGB1LeXnzEgZIpIBswhJRNQdH
71TMQbWnQ4PhOPluNWOQhX2LwpoX1xAfU2qf9WIRCXD9JSDMIKp7YNb4U6/WMCHg0mwLxlKw+3t/
z8sMeRkqutk2dkbSWAYkyQ81yly+KEEXJQBypaqm26mfvjBaKh/9rIgQbxgNuWyk+vUlo4hp+p35
CoOR0OQxaSb3faAo1K0VN4WNyhZzniMns75j2l4QLWlU1cwYBiGMddxyq5I6RPmdO6oU2NGFkP4Y
Oi9tgbF/ydkROTuNiKNivsvcG0kOL+wI4NUKIIVnaGBAX07LLbTwbdb5PQbEbfKelZA/qyizWdt+
qgADEqD9ivb3ZLKzqByqrkw6rFPoavQNLBbHw/Iv6QKsYiK082Zl2ru6i6TJ159dhp2tGz+tdTz4
m/8wDgLknZ0L2nyaheXlyl9OuaKXw4HqqYCKPNPZu/2lGvLSRImnZMWKJQZ/Z3DE8yMpmKEKViAN
obtlRtAmKqRTwhnu2BPwXrUXZp7fWM3USJxmKUqGQMC01Q1dC7MtItZMRK6uTmB5ZNqC37HQVTTr
WsYwgurXKnhyi4NVpuuqohgM0F6gXE1m6dVpCn9WkhSheiWVwDVdOULMeJbG85Fwp0rA9BMz1k9I
DukPITbOYXYLg6ESOMXNULXuI7d5W6MKSjHunDTj9y4prNcamZgprEslerOPcWMc5Rkmw922jepW
XanWFN1uA6owYpwhFAjREx6sUrOLWs6AOFORIlF1Q+KTg//U3vE8AqyYZso6PC1tllORx3VXByZC
ODtnUjIAj6+aaG+OwMfcrG3TFqsl01I+13DTatdlPdfOkqnS0rpYV9jFOMb49oyz/0EqXD/ddne+
O4louRGBUYtFhlQOOxieaMULQDrqhH+ONqdM57/P5rphht7OQCL6tKEyCyVy1CeQ11HdrNHO+lgA
f3buj5JzqPSKZrRRlrdiNOYDFPQzk+/ZU6uwsiA1+LQm99X47SlycG6TY0EAGQi83aaW/JJS/uUv
aLkXhlCVf1zUDl9BtrJLw91uUnmrKhbNNyYDoNtH76p3RhVux8v60H/nrV2/mnves6WQtO7Z8RLS
5FYjbg2bgeA+47pCIllbYrMJJU7TjLyFGE2M0TokhIUXnhhidyo4EATLnL9vFYR0fPSGv/MMSNq6
n6gQDTEf8A8gcP7zvdmHrlxGnp4WVWy13q/WxyEeq/eP786Naw/m7WRIgxZwkyJdmjHJno2dS793
c6r8hLCMbLlQ1Ts/rkEg3UwnHn1DiZ8YnDT8BpsOL3GkS61GfPtRLBuZjGHL2wQe9DkD0mSM6FXh
A8Sc+z1ByDcwppSzbasn89cI0OCJxsco7sdh6m4nCA/JYrRfT70G81xGMLiAAdMMpiZ3UdEvl6hC
rtTtMHOFcaWWxQs9AfEjqknWvh5pILrv3tbpKtf8uAxY86GqgRBSMzjVt0ozSVGCaeZB8nbXbcJa
lqpS+n6w6u1hulasV6zhGWK6elRzUcg2vALHS+ngBDweAT4beXE1CmGIitPxOewF/sdEABShRR+s
vaKw6gh5PQCvlQwG5nOmjGuOyFKeGnXymBMx443fVxdfO1ateu2rPDII4HqdhwkCxz6z3pEG2Mu/
JlwvPnjL1XwwJKoesTVWuS+I2xFs+eRaUSn1rcQsERPAqEbqiX4dsM2AZNOHd8mXjeLn2ZMJvuRc
TPcCbHLw71Qac4Wb9YP5vLlhZNdz8w3TEo0jHkeqn4a9/bEHGUpMAllEqucw9CWSq9cGD0QD23z2
zB1PImrimkr/xGsXe68lK301aWZvybrSjuBCwvk5pznIWUWfojz6nEqFJVWYQV6aqqZ7Z0vAJfkr
RrArMzseCX7JkPo42FBiJGc/Ua1QgGmYEPKJoCzGEawyA61mHUWcE3FMth2O9g2l8JI7KDOPEfCp
m0kvisLPIPtSHADl5IiuwIDxUlShSaX056qOG4uVxIFKqWdvjV30JE9BGyHmgXOqc0cZLuZ4LdVy
udsbDaqOetouhYU/jXkRdsH4Oj+er3NWbrV+nXdBcCiDbjn4zWrALFrT7OcpveqBlBfJDCTqwknP
3JBKAO1WYyquMwNZ5HtHXY5JO3QOu7+MNFgUB+B1pPluiUjPUVLoBszsh2JtoadJTnM2amway3vN
06NAadmjmo84DbbpmOm2sDHhKqGG+rMDowRcoRPjMjShcDJXjzuCvnqoeAuYxEky4EfS4keoS7Re
LOatT4nREJabvY9OzzYXDoyHMSvdQxZKVDza/HOeB7VqF7l/sbo0H5LX7gZB4ewC2fDJsB5Ub25H
SYuITn0GzTz+RUnZcJqPlQszj6G813HEh9VKZh0aMWB06bDoob8UHHGJ5zLBVupieTD68k9cswpr
URjUmvDKj8164ligkJWxMCv9MPNbSxm7/LraUjAaZeXt9CQvgJuaDqgjgxc5F20JVMjRQuiLAy2F
PLmhoyNNu2FI+ycktOTDTASK7rlFI7EJ7ISNXXHYC9VTVUD/cSCaafyRy+263lYWeMs6yKLGHVFR
vHhHNdcnEZvDZuoAtMQCeGfeq2hMpeu1f5m8q4cDWWCYOt3XXLGC4bvgC/eXWcJTUgyVjBcIu93f
UIhuxif5bYiESJqUpN0OoDWUYd7IZxcYATLW6zCAdpXC4TBlCIEy0VtimqX6bz9dYjXoCBx/bZHW
dReB9yFTIVPppageFW+LVE0eeYsCup8ouMepFhJVVm0El58NT1yt7ldj/rUHuWlgkl5hqhE9p1Vl
cad+ir4yMhNRig2Td2E+eWlcJUeNY88tgv/gNdakZD8HwYZ1qkvAMnV900oel+8VxL68kmXojMeK
2oI76rhsVwkquYUNyLzOEcWCq9HnY/Rl5FyRfv3yTCaX57uLSY2L+d2Oxv6Lrs8FRD6UoYbJmHgp
rN3jHqOUbCwIUrO6lVJAvMmh6cnjvl4O3E0/aAydfhWTVWiYpkB0ZNVfV/2z0TaOjLoqlfl/v8gS
Yxk5p2ouaWuCwriVzP5g0KvY1T0VZSMQKtQfYiNeQDl+Q2GCMlhkjONWkD7l3QBork8fwoW6WcQT
dxlxA3Aus4dLfxDWiOhiXIjWrhCt09fVrXmdTHrx6T9W9PY1YFC8zSwwsAbMy5QhKO4+32ibSnFx
5/IICay4vtHi86H6mBVBRZyQVal+MmBENjJcHD03UbZBtMD6+I19QoQNbxRbkyjcVbjf8aJW9S/+
2Yf4s0kLOhUiPirWzT2715T9wpa4bwGM9xx/url1dgXtrJjSCgWNW3kFI8aG/xXuq60PqLAYkQAE
7xK7+Q1F7enzn59aHT2UYG7433WtG/sDKFOBfz6lEK883mloYDgfZyPjtxGUg2KAoTKs+R3GNK/6
PCU6w4EBJl4bPg3Ay1MhIrf8XDOM+y3cNg+W3oaFAxYL0UMnmv0K14rhW+g8pk2L8bEfobwtLVXJ
dWhcvl+m5GGt3KhAASeFVqUSpUVqDidSV4Inx6uAanoS0OrJTrSfyJAUcY6Edt/JAq4Pl4Qp//NW
n3VQtnGjHXqRMxkGtJkqBLqYd9Ks8YJpHzQLbpVxmG5O9n2bKCSmld9POjxIzGeZsUPt7uFvrirc
q9whAk1SnZTYE7eeafegF7pK62EWxNUFEbrYY7zdEoYFvlujARywqpkW2Nxa3c/D/CpFRHN0oxCr
LXuhqlZG11iruT0fswA/kT7LNAE7TJ+IBK3nL4Pv/PL8WQJfmfDp5/PlhoAv5oEyVKV1KbLRT4iL
w3AqhifUPhqHOThSz777XyzKa7WMC6I+n9Yc5CI6hqRm96oux5avLHZTgQDybn64Fc2k7urz7IjR
vaXoEFy39GObRJU4aYM+dhLVzbSZLA+BkPvUWVCQe6qjpmQCDzyKu8bJtfimhRT1doAOnC/YL0bl
WIplA5tVOVEhN3yUKE2MOmnLGbCfl5c6SpFGbSeNMei78qgPf6HT1RH10iVd5ZXlO1C6+AQziyT/
z0xtirBefGM8N1kd6TfkADDff1E42C15mzu90nnQ5s/b3lCrCuJs5ES49HmlT2AZfqnsRkYd032B
pq6jHZWQfWkeYRS1F0obWULlOERaBZXKxDmsvZLNd5EGKaXb9weygAY/z+NsTDfCqJPC8+Amvhu4
sHPwHm03KV7a7/djlqY7kuIkmZ1H53NZWbw9+tmAvYFVz8nx+M7FpKUjc4RZV3EhOqLomKuhhUIf
kMkVOWgiGTKkHx+38phiVPEyHWEZ9SNM7wxHPEsRJJHzvfsxOM4DhfkKtbNUF9jCir6F66rwCYqG
PVGzUMy29XhjNCdpp1deRBd5F0hlZlCBSuFafHl6A3EysTqQ1L2QhLt0YaKnl4gc5mQb+VBTX8iy
0iOKzN/W9TPaqtz42To7cyer+pk35Il0DP31jZkTk6WG0ICFhVv/PMV7eOEXD5iRzoy17Hx2Dlsx
I9xHuzDo/rRAqaAtq00KaNWYaOrvPOS3S3u+7RP2aqAoj3TiT1VogI+TUsYKRBmrcYTOZM+qpX42
UTubEXIgZbIemV7881J8jhzV2qblXrXwN5HwGNEzcRyFqREmHjNSdFBjwIzVFuN5nOFuM6ZFjdys
dsjM34Muw7cGjdlfnrc4oCH+kO8X71ZUPV+G+LDxVCtgk7gAxwhmRgJYwzBaNkup8aFGO7txo/+V
7GKuZE2pa7G2Vtkzh8owUS6JYJOmTDBiYc3+2Qgg+CC52lpp/LtrPAW6eUCt1lnhz1t5hwChlRbN
WB2CkIW5a8nAG92ZTAH6S9nxaFHlGKYupLQ39yf3VM/Hkt7tNNM1ipDIuRyHA3U+IPy2/tAqOior
8VCGzyRNbfJqfbu1cBYjX75JVE9PuNrEPvMUJL+monyxoqW2kmUXrphPJVT2UN/OnIUYabkT+e8L
6mJ9HMHNVLOcB1yYiBxhHk0nhFl8YHu9lhLxTRs3TGTGn9Ey0IgWppM9yv8nTRWNtN5H/C1wmuYe
a//JJgXxOrxpJAdgQFIQOYuCBoRgMBdFGzzYh/FuRBvPi0D3ihA2CVPsLOJBJ62yMbEHu+rRoXIo
cJaperbvu5AQSZw1BxSi4Xmq65+DXUTWb4ZvpJmF57mxEBPmBEM8PofwZgtk23qiG9wuvNpgsFZ+
ggfwwgvowDzw6a2sWTG2tFqpAJAzh7kYRqiYing6a/ditz+DJCY6aG+c7M7dal1cCM8rTRNv4Lt5
B1TwM73X657uUVUgK8QqxJi6uuaDmYV8a7i2tF+4UMFmBfAzF+0QkIXc7EzPY6aWm3Cm2C0Gw3Xz
cBCJ0CeoUbfOs4V0Q6y8dBXtmgnIOkJddHrCKf0Klj/dQtjXujnFRih+Y3zHlgpx/2YnYpt90VKk
HNVnOyxqxIfotLRnvylfdaMP/hrDRPfNM3iqwS1/IGLfeU4jYp4rQQEjxWehrFWQ9lGifnXmR4yW
bqeFw17qrJZFR7nzn0mKqMeBTp9wlQa9NWiFenbhaFuXiDHvdBwyKZu1IXhE4N3fmcusZij0V1bc
ZY+2W2rL7JqSIIkxNjRbH4FDX0opCC6/B9r3UgrZtfO6q4CYbPObsQJS/2qIvzEwupbQx+VOjprK
skAXa/1/ruVdZREib8qefQ9OsATLfIimGNN+HOljLQr8JAK09tNfDi8W76gijD+GZQdVHBTdx1Xy
Eg2chFVnBJV+FQ4dO+WmTd/8PSmAjjOcj53HgdVHu/3zgLRj7URCM2fhxO4ZyJl7iZNo8pK3fbZC
oB6OKAhfWBdjQPsSk2rALnnxZGqabqj5GiDpOZQuqP/yHvtvuTw14XlQy94SwGRJHArj9klZtCzy
/skluOqXNFLbQNjsNdEu6W0f2AngT8wvky4asu76APDZX08mGkB+Qk9yiobVLdXIQYXKURXH53Em
AX3MfaR2zanLhqhAK5jjIpyE6J9ihbnNSRdBtFc7fgW4jwaquwz/uRFFiUVHcK6iLPkeeVfHpXMT
qMjGRl936FC3T5NPGNM54hCFYISATTOAdqKdeM/DIxxomU9Y+VCv8uN68fp60N+0ybqzspNetRa3
mKLK4v38w5idM5EkUudyxijU46GmOG9hJttAuGAJkMjeBDwueibkkJw75mrWcr/LcVapsq3EB9of
fyNY4ImG9l6thpgbs0UFIYTQpZU6FN/UbUSinLZF8ltTB8A0g6BeMa+R2Ez4Qj096tk6sqNFRG9e
FjBRolyMd6f0TXTrUjSi0YwFlxb4HL0EdKYsDDWTXjmYnKivlYpiq6hybx0N2pjEqk4jWJb+gMwE
XPRh2jt4nUFBvsAC2TMadkEyEW/pTJQkW6LvTMaGgpu/g3SOHuHlTuatF8zZSih65wGt3RJi8zTS
IoaWc7RLaFlcLCUGYVZ+i4feGg6sEl/7nYQ1HTQRRrOw2IkXykmoqsW3fJmPb0FPFI1RZ0E1kSJp
An5jnKv9ADDU3ZlnxlJqTT/EtDkLxVD207sGUieJfGbsVWgS3YuEYTNXpGBeq+zkWBRXeuLCdQIe
/C4DVNqe3vPFwKMz9/NWgFMThXhHUUPuewqlaHcyLOxDL1tDMeTUAt0S4tEkiiX70CTzFlNSW4Y7
dxYVSMliqzir7E6cjGWN0hzGKUJXC9OsdDvG59uTOhI1cKs+fEb8VUCqxdzYViMztHwH+ze6OuKz
ldS+Riv+57yUXkfcJZ/7Yqi8hJtxoy9BhLlW8G3afUPQeAvfS/S6BdLTPoBamZvQhvtGQOJVnnKz
8IJ2kS+N6shPs2mS+QM0DrNFBKg0F1ah18PHKVBOZS0coG/NE+ecGVI/Y4y9bSx8YmPmtGsk6/tb
IGwUgQuUyu5Wl2Qw0iZd7oHJq9oyzdckGW0jeb6vv6THf/VDkyRkscok966yuqfGj7oJrf21gmc4
xyPLZehtzydTwSmydvGL1f0Z4IWmJ5Vkgdtc31WjpcrQ6I4S/dq0I1Lg7CWKsOZP5vfZ71bQNoKh
fstoe5IpN7jl78veNIJAbdUzmFVZPC3BIXY4oWjc8Zl1RB5EL5C4hD6OIVYkRZs4fK6x+4kWms14
GES4WfEZBm9/5HlwNs8jDWLXv2KYlElrz1z29p0YDVcUYQxaCeY6Swa5gedSZtG4WsrSkiNajC8h
O2rfWBLukWwHu/coFZjYgQjpe0Bulc3KbM4KxS853uQ7I+zd5o2PhbsYE1n2QZ2nWDEHa4C4zUy5
9dJdDLGalStLGsbBiz8nFtSecLKoq5Az7qwMPdYCbTlh99rf4PK9FpuDyMC2ungerSVnIn7alVsy
ntEkiQWG7ikhghelU0kX/W9abbGGn8DTwldOlBSLOKYSBr3qw6MRQh9UjiGDuYEnwYDCUEaGvLij
GmMjFWG9Z7edOuyvqk5w7OEaeOw5icv9GsAxN3yzvtv3vW6n3vWYqWehFKrTGgOKMuS/MoJPhNi/
KiY+cPwXOzxtImgf5gi5M8oD17gV8N1SrLws6tndaOIE2DiC2B8bcA2YOk/bLol1gK7f0JIJOkxF
jD7ZfUfiCVgkaX8yUAh7dPCTmUu4nuELAbjX+7q6vNBnXGqw28z+nlFKfyh9f9yS+nbjNDKKOGEC
UIalwvjbb5HLW8CKVSZXU3aDBkGiQwgC3S++vxYVTZHLlw/dVJoHfe0ifgxBzBLUm795l2e9mcNm
MOXk8eISiM3YUBMIB1u8GLQay6R3tT9qAoicY6geUiFQer07fCj7yJgF7wjL5QynX0JtNN5eWeSB
okGCuQk2gInlM3wXXosWD6YsFrAj6rmV66j3aXq2nMJfYoF/iOBWAzsk/2k8v5HdAJHN5ZJo3Kst
5y1BVEOe7XSG3gQIr1PiUPUHUKQKzxQi22v+2+s3ar5GGxGAEBVyl0TBLQ8F8nWxijFxpjMHnfx4
4joX8a6/YofKtyWLXjMSQBUOYGjWcthSzlL8NtALVJyeSGLQSJ6yuxcWlqgoruEl+DkSdHTi8UWa
B5fDi+Ia6y/yYEeNEQzPj9FYP7CmZNgE0SJZ7mhYNVbN0qV4gDtn8LEvHBQIaJ8CnpIYxg8tmJ0M
qQGqdCNpNTjCxxokAiixP31m7QCDnTTzPw5DvDAMm3imIhdGwURkTjkanPUVs8TIot1Xz+zYPtvT
nDukUpqGlWCvwnlSoTkdwNVRSaJlqKCe4mRJraZjGQWkS3daxjf5zII4fcZ53HeAVyAhq1pdHpnb
dfyoRWlUS41IGIYcckeFfQOMYjklI/VqN/PKHzF0M1uzE6EkASWBzZtYDh9CJ1JVvlpOHs5mmFPQ
98qmIJ0fmsYWbu5ILv0LKOt+x1+UEN4JALUIFuFIC35cGhzUCccYWKTvRW2uOQlwPj5SIJ7DbvIk
hLfuXkzFlzc3oDEYE0eB70HRM4cysAwcXzw3rcfmk4LUPV8IKpSXQ0pp265LvgNXznaheTh0vt1k
1C7SQz1Rpxel0doXsSy+wPvTd6ZE33chxDsBaFIWwctB95/pk5fln2UKEvAggPmw2BBfSsnHkRkL
hbA2pCjKnZlqg0JN0XRi+58xz5NNZHH4YeLVOJn2jRvMVKK2rHLfTPvCY1wmNkIdhWNy07sE+ksD
CuQaKfYbAiO9MH+hXnuln+AuHxB01RK3Grm3ledWZUWXh8s1IjROP8hut0FY85vWyFV1impKUr+y
j06P09WcSuXRgmTy/cDbz6ggA2t8Y+PI6iAoIjdXw5J3Eu+1vtCKwXbq79U60Mrg6LYAsjUyphLJ
/ppsifLYOhw5V79kO2MWJV/O2qcrUpReNxa+xPufcFSJg8XDAvFe41KblgCHx+eJysFtnmMskXKd
fRTI7dHaZJr80PAAyJizJlzqdaOrphidvPczrlNfMC+19Lyqo5tK5p1HN/tKHqQnfJ+0nvF3lhbJ
AQXOWOsyxTu4Ek33blCxS+Mlb34eBMdNdkP33/U1OvlI6Vjdury90B8QNRPpgPFw2oe9V5BMs+Uu
nxazRkyoi39BxuwrqkwPfpmPI7wDFGapxMHwfdEieRhJpe+bsSI0NOIr1juHQgWMGj/wQOjaQKzH
b8pqPQiZfYq844z6YJQR9i/2vi4YzpX+29wWWk88q/p7P5Pff8tQehXmKXtAO5twHPc+xSNVrYDs
E6ZK4r3Z2/Y2/0fmFqOHxi8NLQtjV9osdjJgL977xPNZvYgktBzekNrr3yXLqZF5MWPIB0Gyj8aG
nBxTNKmY/bgrf1Urdc7tDBlc2z7GCe1pDymqFK8T+bxdZqQYFJdwk2vyGUcmED3pzdrrwF5UM9nS
JxJ5gg/hhJYU/OZZ10KF7fK436NJNIk4t8peAe9EUAUHtFn6+dur1VahdWXpGri3oho3V/yBne99
dtaOI/O36VCJeq2lBD8CjNmnFPIUlck4EJ3VWskleM2G/X3LM/ufII2UebZld0S0ySgO6k/bhzO4
jYefsqU9NyHLzyKpKvyxAudWmxyJRN/RCLI9fEToy9mMAM7xHNlBK1sroNEZPEG0Kq1s8pAVcPCC
YalEM2ESJ9XmRsUvxKgZUsLbjYChfLvk9cRXD4RBis6og4nEJJJME1laCc4pcdRpLqg3vcGYQ0Hk
A7ED/TYDcAIwS7647gjJ+VZbzf8QTU9UhKe01cCdBks2pTczOeYxOxVBYWY6ZIJN81XzMv3KzRL9
bUE4uSSJwyootzuWbNBZBTQm0ex91BDTOiVXPiGdNDv3oKfZ8VFuhkl0G87I0U9Hbs6lUsjFWTh+
yDqayLDRR2KzwU4FKxJ5GaFn68XGIS9Q1QUhlSivjtYAPCD+YHKiEljx/J6kQLtcww9v1qZAYeQt
R5Me4ESRKifJ8lf3VFoC91gFxh00vjFX1oKnNXgpzoiLpOIJS8hyjgtp5ihr5V1ribjX3XNAJXVu
KQjbN6oiEG5oivGzG+kUGH1PY5SsCtO1sUX9d+m17kO5fYsXyU8olsex53eZFWUdZmAcltMhMIci
4lXYTnzkvtpdqfXjD1AAFdaTvzaBy3iJbJtf68Si5yroCtHcZd2XHupycpFK68I4gWBa/vEsI9Bb
Mo3RopKolBpcO+S7KtAbstsWHNzCVCEcreGdy5O7OTGNH9avyKWrDcgYF3NAKcjmg/LMinADIMMm
dV9Rzr2oE4h3WGy3FIp5Pc+rduDgtSMiSwxoE2K+Jlum96ttIraM9fwlMWvroCO11VXWVHzFWn48
FIQJiXOuObnjQkHb6TqWBnPUq6289Uq4Mfst/FENrkVLdUwrYMThktqWFCPm1q4W/OKQWUWG6MuR
EAX2Pos5Qt9HCurwRWnGO9uOzUUKzRNtfvZAmzjG3tU7VFiEzH+ptOq+Z1t9Rbw0jqcEHt8J2Dbh
n7icR91M4yNlL4FfgnCE1JokSnEnqQHo5NXrq8BxvpbHYJrS2vJyA/nVgI9NG02Zfee2S/W3HBuW
j+VwNuMCc8n1hCigmRDUDsjH+585ayxRQwZpXKgbe7gNUYwtLzqddbAQVPBqJwWdvc/wGdUpFP+j
/RILUFqB+TmUcmpX4Yr9LIY9YsNLgXdopS+GK6zKFTX3OZP9aQzWh3AA5NRc5/lqmosCqjnt/E1J
Uf+LY3sCZyTyIixJ44UYgIvpWjzkmiGA08CBdeHp8m0DQKuWmN09wUx0Fis1qTId6BTwN35BqOsJ
u1wr3Jo5StmZFGkbLhUmFkWkGkvB2Jw4PEfcS60Nc4OB5OT63WUR6nmESwGINKQIpwMV/CAacXhj
qBqviZV0jXOABmE4v8BIQ+S5M9S+WQhKN2PemXZym+l2nsS40ZdLJg+jfNCtITj9C6gE2X8SK+eC
93UsL0ZPYSr5h85VflBvnnGkYyCCuGe6Q+X+mTf9qk0o0pcIkw7EvtrQlJcULQ8Us2dy5EVkmDh5
dIqZcmSNGFCC0z/4t0PEuOOJas4ty/v1WGR/2fLoZ34vwYWT5R06dyooHTCTCbmIfvxUgVt4Zokt
4XQMwU2q4u5FahCDV0QSUcJmimD2yttgBd2/NrtFKp5O/nGXkV/57pho5aaLkMJzjJ76/ZphoNxr
da0NJ/7P+RAwWqOAWnZyPQ/LXRQYi9wvRsTP1cgBPZt9yrzs+wqQXtA/LA2Fkc+zGaT9S2Xsbgwe
oAZoLnfQPK+sB58DF6uao3qmwoFezA4zYFG6AMUNCdgSCy9xUuCZ65zNWlpRHHpRceNcLe+HK5Qe
rbIxlMApKn4QxfolMw9PdRyv24ZWdtcM2H3fK32MJnl1CzpxrsT6spNIUW6b/wbdvwX4E+WlDAEk
pRAik4qPUmxILR8bdJQ8Jpp1kBQDS5uEudwg0gPmBZ3Loimmi3l0CBflfGvrPoE0PFkejPwMxovK
ZU8v8Fc0bnDU3UZTbw5SwYv8tVvEb5rZnrMf3EgaxVmEg6MFbIXudowdfZN8OcdPEyuVazwVfn9q
Jt6PCocCVw5a7WazVetIHpAYHcxT1eUipCM5wURwdd2diWx5/vfKhMz4m1y991ZsxI0CcHyVDv14
tZa9CiisFO7PNJAs1ooYPCS3AnS/aWz7ujP8wmp0EvaTSKv4li6EiB9h/FfN/bQNxGSOtlg5YY4y
dgdYrenp3R0sbFwM2jsgaiUTjNe5FPyT45drQwI8Y0lZfIQhzE2Ecl9g4M56xthFaT45p9sQmbTX
qD89rapCTNQl6zhSLL03nLJXoIoiolyTUCt+VFBtgTBcmhdOi4q3FsUzDaU0VzxOBrbjJxYfWrvr
dAkLWIGVk0IAmhjsWUyQ8CRoKJRo2vNtEKad5vA/HK0tozQpnpBkR7Pgo/z9Tzpk/Vz+FgZDp026
CXFfUo+Kmn6Da6+WTRt21aeDj9hWJm0ogNK/HiiIx+BtCmSMTIDT7Q7rTvYHiujzWwMp/SDxRNNh
vqJbvwQLuzxcZpOhEWyiAWInxSN9u7uchRsOFBXcHi8ysYUqF/R50ypGEUB9lVYL0wz6N1VGAeQS
Krwisb01AUy0+WJ2GHGzoDLull1b2y+lrw0wro7fkfk3bB9JBiqVuxglBNEgUO9lHMcO4Zd9LM2O
T7NcQZf9Ffw9S4xpWZSHo+UqU6h/5BH6ARkKtu/l9NIaIsTRyc2/owIyGJad4uEiAJO91jLxqE4G
YqU7OSJ8SkRXLV83MKf2RT0eUDrESJLU7cK+AP9FY8aQ/32tAe4p87nYO9IbRWkhi7AuH8PBKD9z
o9MvPy18IFsDoRZSVGh1OVbillq9AOdOlT4UoYqlALtUKEE3zsiqPTr2NeEOlMrUuGpqQVbQHXhb
yICeYcLlFPBOSVCceOu7PdFwdH4DHN6vvgCkooQyAtXystFYI4zTZYhXJWb4tsgExLOkZOGlVUzL
sEqA3H7N7KN6UmmTiT+nAwiuZ28h9/4v8tpkpNMOMV10VIU74nmsh5ZMW03mEy83v7J8kSfBX/UV
p1dg1p2FLsuFjJKTOaskO5mALKLf9zfdABMurfUnkZOHvZu+sFKn98LwurZZn95TdAt38VEyGj/2
PiQL0IOMXTN4ZAQY0KbDxvSch0RH4vxZq1nyqw7v1xe6oTuZZ1AWzkderLU3zNIjXnFoOszWyoAm
lpXisZbVTzGvultEIJBNOrQ+SJR4yxDVdwBPvU6aQsFjVeE60FsV3LslGzm3C/i/wySZQqXglGrR
2jtQJ4PXiH8uKCXz9c3SsQV57uXtPvx4u6bvjr2PUW20NmsFoSXSoNqlTgUqs2bJaaAudXj2A9tE
GbFywKZbYJYK7Nx71TE/LJYhsV5CRJ4Eh5IOaGMjETkEf9OapX5juxJTk+O415gtPiwYEYNA0Dcr
BL/7Zuhwjbuajw767bTnfCazcOJnIeZzjstGF1fwJrdBqbLbc52e3bwX9kKUIUIuwU+cXeQZGke4
jsNkKw0PdYxQceC/SEaeafGq3SJAUKcddMxerS/xJ6LTyQqf4XWFoLH44pP17hdB5oN1RrLUfwOr
6BcXJGf03YCgblAAhMd+Sm7S5uEuY0B2SJIIQ/1mLn7nPUCzRZuPl0a1ZX1NsNNaOr7hTuzW1ogJ
oK653SrZKNdqGqQNIyoqhh0t18G50abvzR2bJMIKbLaDql/nwUQYt7bwCqvQORjF8RW7JcvtayG+
I5IVPfkXNvJmPuU3znnh4wvuP5oTrNLAODxb0oikYA1oBkqWbvucdjbvPmrpFQfdXswt4H9JDW9u
vpcaBEMV5WgQuM/NVjAAQWGljxFZmXe+AAjKXtN+1d79iIP0LizZPdDYrVNXdxCL2bOXCXz14PkR
cNYfiMjv4H7gfmdHHBEXmzzTCX72602hSXjsKNXfnKYx7RgqE6AIgKucM6966/RiPt3cRnz0xscd
dT28FvOjP6GVvn/Tb6SN4+D0/GqP6W1LMOFGKPN3K8r4ZEuT+DvqifF7Qfg2wSLL7/XQVnrwGARl
GoSEpHz+tS2CIk8jZpsH+Sxto/Cd1PG+5jRJTUemQa0/IVesF46cShwdYaqPLL0F7OcfnbeLWu6Y
/pwmQd8a/zryJnxoPUZTBqv0BCDYs1kgzH7jwfQkhHitaesqOy/Kd251rMwEMZ+WsI1fLfUHWNdL
Wwr0Uxk1pVSivk4Q/20p7UqxYBCuMroOvvODhBqRROoF8/3cS4p2LutrMzp4ZGiYfwXpBxsT1xrm
MKRTvOchyddp3/G1EzAglSHuz/T+bEmFquDSEXGc6ZQv4qIriBMNTn3zQMa833F139Wf2Q5yqVF1
qmxm3i1ACfyzq5Zq0wIKekadDYWg2E7lqp9YaxYbj7QGH0AMCsSXLTIu62eQ1BNDd0H0dqhZIyUy
bjOkBzTXUoFEDCO8NLWFczmDdbsXIp6ccN0bEC51vBZWO1YBF5vxA3IjoqClYibnpJz5mhRmvp9O
qYGkh8xXpTmuRH7Glf7WF9DcnUFtJgNeFyoBwamv5IVcdvldGYasACCia8XHhp4qUKM5kd52YKtD
Tt0J+VKEdQ+knFBmCEsMJmBoZlf4JrdtQ79iTmJgBECjY61auhIy7Vw2O4UkUl73rlV0y+Kr0wWL
Bfh4OszGZhNLtjSAqdKYfrqxsuzsQX5vIiQdTlXVx7pjjwJeozRbKt1uBNFzgRs9vefhNacQaVau
sWrumaaH9wYB09Wcg+5NyeixjhgQiJgT7jI2tMlMDJ/KEN4VPg9yUkJ7PC21cE6BuoW9PzO/ebWL
Rf4bxooLqlaShglB9YJXV7yoOelgf32TFZQzPW7uvO86ATiXDCGFqGFGVpXAnhBHXGbV0vK2Wrup
1fI2PDVviTsbUn99UYhIuIQCsPAZ7xxX5GbG9CE9IOjuKjU1LqNc5TyaWxdfq5r8KoHXNWhy6aS3
br0yh76NHGzB4AylbXHPPCGUoPPSrZ8eP9MKTCvE/i9TvWLPyh9A5WImhyjBE3mRIBenOjqehhT+
nnZho08bOP2FEXK5eQlS2t4iyno9P8kyNnEihKj/Ul5U+wCbRSz39vpdk9TxzBm0UAPD0gUcv7NH
49orXdEjHaOhhqeRZFd57jMnginO2pbZrABD6UlvH9OUaaHgtazx1eOh1WXR8S/TEt97ky/dQzMQ
ne+EWd5WAKi5V1B7jWytakmQ8RXCugLMatMlyLCHxWMikDjOYpKm4a6X2sFtosew6gdob6cEeDaF
WEni9lXtVk+mO2CM9Nu46hFJwl+n//NzqImNQyRd6Kr/r+sGr7fkBzx7VyKnfPKdr5dBXMDjIM3a
rz4OCp3bIrNJH1qKGZOicKdWomIepOHWz4/HTwsSjoKCF4wQqufbtMvWGkF0oPfMtLycYgd7zDGn
8fnX0hsuvb2XmSKKpVtzLyUklHJ0fm7c3IPEmZRFFtL6LdV4380VOOhV3CfQ+eZfMeSkf0M42QsN
UVBwC8tTOsacNN7z/pbzeUIit2ngNFC1h+P73X5OpvfuLZOsXt/dvFfMZ3/plGi/EcXb6MxUC3/z
0ywA/0zC9iyJdwxcTMS1fshkH4DibCWPKtwid4TO6HMFtdvOJABpEMmoAhjnwIWHIAuEeV6db3Ve
PqEGS1150CocK0AJrWl53xVF7Tzthodma2FEjnopGZWS08VPhiP0bsj69yM2hFmUfDYsxfzCGkih
0uHJFuM0UBpNMvh314qMHq6oQ6h2z7i76ic6Y7zJoAASsZISsTDGbVaks1bZBQPuoW0YyImZwDpz
4xCCCrZp/mdlvWaUMA/sLcRJ2POWxTom+bjWd4G3reQDsXl/67ID2IIOq+8T61JwchU6XQy54vUz
41BbILSeRrwV1FmswV2YdAfvMTJI8J++MlxpCayRhz8X5gbHCNCKEN1z4AUatnOZ5+mWhVRAoSwc
h++s99fSEJADUrvyhp3+Siph3NOPcu/20rU3VCChRWBaWGCEpWpN/gQFqedTF/Ix6uYRVdm1iAs6
fWSRLx7wdYezFEfsoC50A8uyFs1THFxLQamfVFYRqiAmTCOg7YTHiHldVHdUZW03lZgRVk/wAmQn
QO1G/Jqj4NY8GFtpyePohkQdO0pMmc3rrXfk3Y1+95c22rA1+ASKjyDidPjOmvPqWljlsU/5lj5E
VxDdSLYoLqfsBlSnXiOA8qEnX0ieu8z53pBeAl+UU38M5G05rABomRAr2dvkHa/0ra6z0L49AMtK
FGx5WqtepbJz0Fi+8kzMrp1EQEsE0qzUoowzzC/fNJ2xADJ1cTQ3eyL6B/D7DnYqtx5NaCAwI6P5
ZLe1k1QN2r+QvZEL2PaUhOxDmwwrLq99qQ7CeT6mGlcirpHvQt+i1g8f1NGVyBSsEfOOtStNMwBx
BUHX4OTRRxNGvz/gtT6WWvmotOoEysC49d1lHBmEMxij4ZtzbQ43hXjmb9ecjq7oBXMH+XfIF2p8
xaYBcZII6zZhI5olaOsTHaQWtQNzfkUDbWfAv+uQgenjJEyGZZt5ztJT+8joJzkpzaDy1DiI2AGv
HgjEF4IEEBcJll0xfMjImLYrS2VI8xj0aWYytwvm68O3x2sd1jSf+AFqj223A6r5X0hiuwLBu276
ZC2DNX1MzNfSY0UqfbIlQrRQPLbopkcNLiVmGkVC/+FdsqglftGA5TjNS9pGOrcWf6rNmY120A72
UnmpG3qAkl+flAl9C7/84sCfV4ZieNowrYXeaQVPU+3yPjk2Uzh0dcZXv2Nl8JhAXb17MrEuMZAr
q9dvw65dUGfEUcHGZhPa8Pv79WurB8zVTeTJYm1GK2sw3qD8qOHHfRJQ3T2JOzOyox/mVVpfxltP
3EAAYk7+CNRrkV9xbvAf1zzt2mOZsuU2p5zhNklH8lI9cyTvuWaDd3XszeGNyPcOMnu2u51F6Hy+
26UEHWy4vQemtsD1Asnwa+4TuTCcRMe7J1Y85y46Y0gWPMvKCGoF75jSSJlQpRF8aWDJ3x5r64uV
+HqCxQrOGCtQBAILTZsfMOyYRUdxC7O0s7+7hz6woknL+Cw3q8LuqR6mr/GXPZevCxkhdcZ7T7l7
oGG8q+UFUN652D9m349PAr3XDwQ8IVEpZG3BZYS2OOCtlVlMS09efTvmPhlyrd/KjHmJ4eooeEtY
jFx+VEbewUlXK+rh5gclKaQydLx5XHFtq0Lf2CKKBT8eV8exF1VszhH67Aw85u5JSkU2nrv4WPVQ
Iqx72GewQveyiRjk9NSBVhNLvIc3gsnF8NywAUrXQNfH4hbQ+5jY99T3+wg2K5wDfCUanxmEAlWy
+inMMfNOx8I7ZUaqgGDrBij4er7hPbREDccWinsooULghMAQQRFrZycOPLMEJ4YJp+6/zKBNlDNW
A0lj+EgHZvEUZyYksAD1L5u0khfL9IFWkFh78kiV02c0KlOBpS8CFKLScexqEwBmTqam0gaGo1lq
kELKmwjt9XpDj9JbWq31PI3wziTM0SeWir/6ODLo6NqpiJqQck9ByS+buf0uhLpJ4AcmK4Jj4Ktg
GLTc4pY/5Q5APIbvFI9mfyNDrw3YRCevIVMwwGjL6cvcbFTgmwlAMrRnSbwqGV9LAcdSuBsIYUGs
MRahjkOAfloiozhzJXm4uexFbBHF4CNpxbJ5ciuCf1noFNtjpZe6WULJfq1RPxMmDkLgXN0g0yWT
Z/tOncZdk/AlNT8yfpsI49KDX96VNTYiPokMtBtEVU1I10NamFM9IodIZaMZZJUvCT/k+A32V5H6
GT7VhWoRQM5aMY4UAcD6b8SZb8C04Bfi9T59VPCPQjP1poR1pzoRM3nZgmhA8cka6WL/R13h7IUt
j0zbQiSeiqOk7KzpD45UqNSz+t/GkgLjxAiOOEoBORX2iLTLeEa/+YQZOuQrDNppGrwq37cQ4Jf/
hTJcKlar2DClxe4vfi+roXY/RDuLIzjOJZhXi1mPAzMzDObrlNnXmNfnJxGITshXhHRapirPiVbn
1EQrtqEuitV+vV7JlCb6Um3aTfU22pZ7LcDlKgSPHjOUq1+8gZpAfRda4BANnuOmUx9E8sAskmn+
Q7lYGfqp1FmtgXdLejdHypBDIc+DHJDzmHXbePpjTvY0sDHEr4r+t8vU6YFe3zmWVmK1BMoje/io
qucdnZI+jm1brDbRdfwmna+Wuq4j5H5xa9CNIF/fskknLpmy9YHpEKIPu9mLVvqCD3SIjbk6mccb
yyq6EYOF2H9LmoH/1bHWoWPZX/cJlS1fJEJxPJZPoODuOTxrXr3RWuxMMitxMvCot1KbxDJtqIH8
+pcgoN2Mrp9cnprJt4dWukHvlyOPitGQHwH15x6CI0TYzqDIIe8YzY12DdvNCE7L6HAltuUtJu+H
fnpadJCpLMf66ioquB1gPzLGt58KLteWaVeNvChnIlnVFt8/XQ7BfKkiWl/sPXVtDlzIdKWV7gEy
KXBiZ0XqIDITG5PROwBsRzm3X7dEMs9HVWGZvSkSSBDcd9WG+ij/MHi1yvRgeS55VsVbbxH8zo57
MvHLdkzGQTBd6FJcBxmCWvNbeRJC0TKMufCWKSjO6hiK2A9pjRmvTNFryWrslGB8oRwsMznwzM1U
rXw+OHoiVt+moYCFcDMBwhH1N1smMsgVAqLk4aZzwMyQRguBnbTvxHjz0ueqxdHlvTv0S6UtfSpa
htY19q4GOJGPxED609xB8FB5+8qivmowARnnwOzJn0pAJZ+tK+lF/7vxHXlae3QR7W11iYl+HUId
L/lEGpZucHUABy4Ny9a+m/EGDKMy/qk2eeaD8aJjhX4R9LGOVKbPihPluc5/BkmtFNg70xmrjUQe
iQpAHveR4/J65XJnEfutbIlZeleM6mn5j92A1iRBsKH+2+tryEr1eBIyRNuhXBn4hUb3quLWfVKi
T6tvlODRYksDHFQYmut4o4qzMxdRM6RDpWbj/icamzcO0nfXw++yJeXTez3169DqbQodolYlrkd2
p4q6y1z6dQgTweWeimSQ52OKak5h9LrYgYMx1CBWIuPgSeWRoMPStmcTp9kEMbXvcjtXEbp9C6gv
tfkUTPGhAZ29XjFqP/Ed7/xT+8OpzoCarvrCsdbae9HpdK5fXSr1GcjFaady0bzMCDH4L5HYJ745
dDT0oqAi3qoWqfEhseU1FbarqhWGV73Bl/1N5bZc4wP9ounRDCvXgmvR65k9GMjyATxsFcWdw/4M
Omgw5Q6AX5DgVBTaucXe7wAxQueSEGK0brEADHsQOTUvZpEKP+6cwPEMHJtZvcL+DlDp1CC2QpVb
+75Bo2y50duUzWiu5A7BJ3Ag5ktGy3E9SvuIFWjAeghSOXvtu7PzqyQ/+5QVqbtzxw/xY9QiycWs
8FhTYOeUdbKAFEQdwB6llXTHfRhULYOzcEERsM24IXRSUi2yIe0sNrhrX0tR8M++TXkRNdVjozUO
dxcxSjF/KNEY8yFVy5XgnVP2AxkDJLSc0PIiZSxV95ZTPs8To+IldHgWHim7bGF320z4apTpquzY
VFkE8PmQb0a3Pt3x69t8IIs8Jmowd4VuIbOqBn5A4vyf18nyQWvxtxIIJlgwVKQ4mkFc5vuavUAu
7K4ozEqbCEJCfGVsL7qPcgh2rKxxCp+RvIqk3piPDRRTbMDDXECidcF7hp4jRivnCm7uz8pGbvaP
9AIty+VPzJc7A7GVXWtc/AbxIHUaX0SDliOI2em7LYpbHTF/rhIdaHWFnpugOTYWSpywI/PaIFE+
rx5LbCCZxUCl9NzToyMvorswR+Lk3tR2p8w0jGRaXhJn6g576h4eUZyVC3xuNgPl5kosuerX6v3+
ACGl57tynv+AFBfm2CakSMkpaqnL1tNHMdQXHXF8rRElYq+SdBl+8WP6Dfa5BVGtiWF5HtFaAY4u
x4knvwRnXcMeRsDw23KbZhEJPnl7w1UOURT6hAdAVJro2PlqelE8nbCDpg58ZtVw7aeK5v89sVzf
dhMIhOqK8iFKWclHs31/DKH8dC/hKsefK/+kB9wfZVYHPkuLcZ+TGQGO+uNZOKOWIJwX4ZgcQNmo
Y2avV4aFYsWt1zi0Lqged6DeLozH5t5zXc1bCA1LONqg5dWPCv07ovKJDQAftvkwlFuyGSIFPasa
kElViigRukU62YU3DQUfYb8obKyit4rKqBWE1drsOfQzKvdlJJXOnukKhBek7VVStLtAD76K3Rur
tsC4/PFswnDTxYaM3M08zpg5L65nTg8uaAZ6kZGNJM7Sqys7cErT4bzOfNV8TouopHcYprloy8pP
jvpUp6C0HKJd8pNNmpJLg6uoWvcPIwfMEioPoHXB04mQCHkI83SKtjllSTKCdNfHHfFx1umHXGjo
xrEVpNBhaWJjr+iRZkZGcU7+ySS8kMdY/A7GfM3wnsV0AYdhyao/dfNTGeq/OEJJmsws4Z9Dj0Yn
We/PCeG3ejP6v3TE6AhLt3CjEOAwjOsmWUXzkECP91d/nedxNrZoRJ67jDZsG/QrfonBr1ogmkFJ
Chsz7ii+Y3a2dE5VYsYl5kK0yF34f/RpWsjKNGDGAE5dtcfix/ecuyHuLq3v2PW5e47uLN5179oC
QBFxjOSHgPG3l/hUfWT/lA7/uVcZnuLgcOj5SxdRFbREXgJRgEokzIw6blUD7wr4D4KanPJdEWJs
iHpu2Ijqb6ucvrTxyWAKC7OAvoQ9/GgWLqIjC8xIgWyksQmHBUFUY2zztnGbCIcax5ufQW8GInaj
8nqy0me2VzeVI/KKSzB+9simCLdOVCFyithfHTd1MznV99DRX3ZGqSRyPByMAjEHgvkvHPOaOgky
Rk95DZPiIYwYMeQDGHFU4r1xQ+PLkBxWRXLmOCZ6z0NSB6B3+fk43rhTjnfr1voS1vbLK9lRM/OY
amtRtmStkGEdKyAaTCZ/2C2eptHrA3NGZxmPYZd2QoVovwCM0JGTmWwF4K2AvnvwKCPVbrsFm8Gv
5gpdJHYyt0ZJAQNxq1z4TUUQCacCJDhKRGsk9/ty6mSKKwr7SjDUXWup6rzndbbjXxmMIcj9jW3X
+1VJefFw1OFjflemSxgWFcbratiPe9JEd5TdVsMliUOQHgNRB69Vlf118Ydff6fgp2XKoZaTBHoh
lL/h+F3lL8dfxZnGhc0XECrK52rtJGOf4uosGwcoRxdVeVfj3tCt7F4ayB7RRjol6o7JTil2k+Nu
/XX1VUh9iEXqgmAlNf0UC7OIV5EGYNX5CPWpYl5cr0hpdbEbv00arTIvodzM1BpFkShyGHsHwAqJ
KIv9ubSOmIt2RjYCAthGqdDdiyudgreamE7Dlhkf62tyHo5qArmG8DvoeRotd1CxEX24mGx1MsLp
SvRQsKj3/mFg1fBnfnfjZo9V1xoRcSTxlbfxVCKQHcS8JvWYYhwO5KEHSRJat3thjbXM9oCFQiCV
Ei8EzT+ZPJhFvMN8eNSAqMYlSNAQDVwI0orU8jUj4w4McJJeQdKG2hvH/xsZ5YYJKzlUyY63AAnz
UmWSoQYnwEG3NE+8caGzC1IxtE/wAJ30kuSKpxT1lnAeCfcS/bT8WJgHRgADPn6ANtFXVH0DvxmZ
iuBscjMx7wfmgVcrWvOkk5oeiDVlj16xISo+1clMWpiiR2Hc1PPnqOOB+NJ5p+Rq744iNXEcJGB6
GoY+/FQxBJQJUhRbBSzYpmq/XxbHf6BHZLpFcLTyFsCIMdIyD3YGZd2tKRuVYUfDeIcOIkF21H6f
6VtUcA+ggAy/kOAPgx0O2UWOTJtv6mFftfKLp6p2D0h+7OOyBohYlx03cksPY3r4EADt3wCzhkbt
fQ3yoQfIs1wt0WSOKsr5et+Y5TgIL54e7iYwx6m8JkF6+vTysF5jBFtUfs31ImIHXlY8jwPtipAY
9arKXdLJxoBb5ni6WUzCRmHsAaCs0Anm80xZGgEgy9/hghQSFbQXM8vR7xRrYwYFjeGg+oQaizkw
CFV9Jbd+wXYURhGHaeajGeesvqiNLTjvmKt0c0k9Dth34S4akdVH6M26awfdaR26MUZVcrxg1ggW
j08gxrV3nbHmgRtMCGDVpp1xb3CLp7GXkZfiV2TyC0QeDj2uYD0L1AtNAMjFEqIHsAgjUrYAodVJ
l5ceXkVwj9yP50y0UOfmvXkfHUChJfa+xnR5CZLAERxgorrTHu7DavRHxku+DXiWRbkwJdCkio+l
50Qzx5MjFzRKxQA2NPAKLbBPFmDvvRiM7dVRjtUk6XzNMVoF9Rm3F8VdKUjfb03PCqs3sONYlio1
dQbztw6/WZGbq6F7SzBB8JL/UU3ANuh08kqg0Xw79uTBP/qX9oMled8dqG+NQFM5bW1h9mIxk0CI
r6iC5BbRTWDXwvBRci6aUDnNa7gW23ND8Kp1zpo3yn54FLu3UHZHtx+6eUCPU8ukwqhMNPD5eKnh
RdLb9ZEC2ffe6dtILixHfxvm01VKecgrUyvkmXctGapssXKu8iTj5IB/EpQwKryHiCsw/gbOUqWw
wR+NnpMWZzd2BRVh24aDg6Hc3PhTieRPwIr/tcmuaM2JLQPAeZwDf5p4qOXl7J0YrIR8iqt27XVf
ZcZwG7PeLuLIPSTydrL4Xgiiq2hsRZUSuoy9xkinh7Hqr11edOz1OsXjU0dV4HnYPQ+ITAu6XKN1
yNf9XknmL1Ffu5pp5SA4LDuLlg1tIlOb8FbI/JEMgQ4F2v6zBeHRdHQYDCzOmS1b6lOGpf8AScih
Ap6XvOC3o8n7zUUtldPAfNR3TFuhWCCgf69bD5eqGMxcPK9VSoUWL9OFRLWJ9Sn1NOXrJgu8qEtI
e81H8Ru2zB9rhSp8BdBuMYVWVdhkfZuAhxTljygN0tLTKUlnC3gCS0XfoYh4WvQ+dVYHHfhguzbO
G/F/em3DuQyq9bqDWPiPm/2PDFIlYqNNsz6uZKVA6n3vk/0VHTrek00myZk949n+/vAPTzwP7F1h
1CNQwi8EqUC+oK3T60maAvMpdoK6dc+vk0D8T6PMUw5Xszd1/SEeNJsbv65Y9Nz3IxTxY31oYwpW
y/KMcEF1aOVzc4F66rkgudEbBy5kqI1lqL6PcXGld/GsVUT2L4rVFkzHi/9I7BJfLmQ223s4WHeD
Ge7zcpZuhAaXT2veNfuEQOYJ2qRcKFFIjz5kgey+f0i39iLdFWYtUuaQh4EQBGHoK0Z+6AzuPDY6
TTXGj5C4Qd/dndvBVBeFtDyWHgnzDIPZeUxhZWRfMRYrj+MrL2UU5CcY/fw+ky+Gvq8K3gyFI6n0
07AjdK+1fzs/obZ01her4myC23cqNDzDIxjFs1akzCP9DUQbnC8SF0WwxbvW2qqGy0ybj1WHGy5W
sfCqMh6DBp2Wk2KpIaJ10kS3hTApLTcBXvqiYgenh+3EDbV5KFMwHrrPGfa7PvMTDS9zTqoPOaZe
jisIsfpWjhKvuI7J28PoDyJaNc9AW97XHPzq9DyiNCtruL/UXGT8JyEp/qct4s5ENZebaWSpYXIM
sLllSeY8hNWNqtcL8SDi949GFPzKac0TEDN5iGNZg7BjBsr9fb3Daov2z9x8kPXjfFiJmH4UGLDF
Q4RuVmZwbJFySN9bfe7kOY6w9vug1uFU/7Wc1X2CJ4IkW3BEFuhUSH7pnUlJmikOYMrrDkfPZhAY
tZVCgOgtUkGCOX2n5Tnp9RHaX0qsdydLsB/Zo4Q0gpi2XFRGfKPNVfGnnc37VgXqXR1M+JpkaIBB
z1LYI6w+bSdloB3wmpL4C7v01hPFs4fkpU7srGf/IqkS4sT5fgolgtBo+XIU3DnLbnWdZoV7tfbE
jZwYC6f9Kri2sdwZC+SCYPMaq8OPrN3mIl9zQWCziQtKJfPyunbzM4b1e6h3J1JiUuCSL4vEYymV
CmyGTzzVz8PRBVXcAHilEDfviULdpiwDs6F0Q/quE/BjLETD1T5dJslr+Che8cSftMG2MH8KeUhB
i2LS67DxoSLjZqewLG5tE/zcfzSVfpsRzn3V06p4KCrECLMa7BX0PA4IGB3aSkm7IJjk1JmSxi/V
v4+w2tWlIBUmOBTisV156eWwVSBZVxeEpH0V5YyJ3PpGRqXBV21VUEdrk9vCSIdhL/3BwDAUky1I
JIPbkLFxGcQpBAhLGma+UBxS8BzUsH3fXcRm1JzOP5UmIbCe2ZO9ZQXASsVeBKGng6e1k6ca45po
tffiYwCNXD8C7gPlXQA6ZDehgBXaiLN89goWrRNi8fMz/A4ndinZNfBjAPwuE8tRmdRFR185c4ED
CO4wdHerrxAl1cBsAqGna3l8hxY+Qhh0uhAgMa+7nEgqm0GRtkOLxgM3eqwiCTtp4x02Vai2Gt4w
otb3IfjHT5/645AV0hepHlLBk3DhADoqRRX/y2p+5q9hFXwKw8MtFJud7O5xAWuWW2acVObZgCs1
FIgmjwVlbw8hmlSiw6VyqM5YAPfcIdwwMWzIeaB60KYo+apMTmjTlwRADj5Q3R5OQd5tyrdhB4WO
7wBSlOuTIKIjiFgKhDwziNXcw9vIjCW+K6DR+GVnGgadfeFUARk5eTBDaEJo9SDiwVTsWwzON2Dp
HJvlhTD5T/5pJkxT96gxpzEEZbvvXH1U2+OCgB5e7yQsBQn4YbG/u+52puDGdF0MfrsGlLjSGvr6
E908Hl1Riq4m8MWHvNtMmBvM+PSr95AuFnVhe/5z4ZfvkUOCiy4RiismmDzT/cR31+nyXhzTDtlz
mU7uXbVzRKs+q1wNidAOk0zSbzyIEA9D55n0CqeCuD6n4OTrGtyldbJHQC3WrT/bPZqyI1pwj7Ym
kYdN3wM15sXkxOQ5TAeP5BUHU+J+y1o8VkozfFfVqT54NzUPW/RQrK5efg5Gg8AmGPjJI8uA4rI/
Ol6uQ1QBbtGcMHOj9cSkVCYoy0eFXGeWiBlAIf7OH4/jW3ASQLg9wp8SoMrvjw7ImLeLiYqi9MeK
MWREecXulX1GFKQiLcTMmItQC2mGc7PHV1FgUSa6Lfw+lNjUNtgCdcq4AryetQhppRl6DAcuUjxQ
3AFA7mGoc0ogYMCeUlR/PH99sAwk0aCTBt9ekuMo1dKSJWHGLMCbJqmkBmXI3HlcCF4hK2JIQTre
IRah6978me3pXGuwQ5l/b627LQzkjW0zTe23iK+/tiQ69OKEAXfW1Z575QTd/eTTGVs3hJ1Cmggy
Ecuh7rve0YW1s1cXp2m/O/bmGoMyV6vvab54ikIuvQ+o1B1csdTWn5iWbXJbKsUmv4vZI07aWU+5
LW5jBZg5GYPTxNaQDcKFJEnLn38gc4nzIl6vYsDBvfzid6fc5fF9BMTGXraOy3jlHSNCJJpOjSkH
p59+3saWPG9q9H6enF6MvIY13kp/TnweGAIKKIc1EirMokEtjS/GB8asPPI156eR2/L6EvtWQrqW
r7FxO6eKoOei5TCDI4h/2kGHOHXo9BOr1l0blTs6YV9n6aiV7DB4Vlxuh2EINGKq1h0y+8ZnfXl8
an1XBnWv2Ni1qP3SEcyZD/fJ09tBYcc9FHM/74xhnZVl+fxvAf3V+PoCpMEVDjxL8jzRmkdklr4N
MTF9UVDIs/FYah+QEhlazN8IAyePTW7LLd5fiDzcTBD4p6g10DcCkeB0sCas6O4QZcp6bPO/rx36
RVq9+LqU5bm9HW6sdeXNB0ei5BH7D1zE2uN44t7GwX9jJylVh+7OwCeWbOvEVoII5eoc2z3ZvsZc
v9TUBiBijKRtIzr97vdXS8fkizWCAykM08WUbEmlJjW23+H0ESGfnWdESXnzZ0UuqX8ey1+y4LaX
pky1qQFpk0J/xolEyApcbY1QXcFsxSuqCClbBNGa3ls8jTTGIRrvDNbEeyOfSg3z4W3T8d2d7q/T
6THmJJQfNqsyc15ky1rMX6MG3Xewig3mjWwDs9DZPCH13dlHXNVvzMw435VZYhfJSK7DMHHd7eZD
b7WeIgIe2D6nC25njYK66ZaJogeZfPV4D9bpyEcT634LAVrwAc1t4F0+ZDaxTog9x3W5Kjn6eOF3
yIkv4pcTchWx0+BuZEvgjx/QLhITTSlKXfauz6F9E5NjpsR3eQpm0yqNAyUcey/LWpXAqfFe9SSj
RcFWeG80YEMiUGlEx8vQOresQxB1NqqF6nevLFj55l0NeGQeKSJeojClP6tY0cgipwNhfr8PfgyP
SoYzHYbzYgzJrlMpGWGd2vrxKThJHtDivyHD0V+jelVz6XPyItRKIJKViGCaX8od1ccSEXBIHjEY
0bwYI2CLpfB1ecTLYw0BWYg7aQ1loZH/yD+zMQqAlNiK4jGhxH+Nn7sNnUcdcPBRhiDxP9nRCZ3Y
WHaE/UqwhD6Mk75vdAvtpj2TZxgJzA9Y6XBpgJww8xZgxv+OdrN4RqunQkFsXJEmMd+7AV0yOw+Z
KHoNYr4TtJCQ/HZgUMft8M9ooUJcRzbNCDxKeQvJmfWR/l3La5qSL0mr9nDlV+9uy67nXqjCemy0
BtrsTz6ZpjqFeIxnmn3bPic4A6P35ZZknfxEObw/jyIF711Ql9KKj9Q9g0IC4gxT09qOOa3eio+E
vV7I5Iq2Um+XawQOVFhseAYA5C1WozizOCWeyBoRZ8xxtBcU1Ptlq7/nut+7Z7d4vA0tFq0yLCVY
0O0zFDTfgpBiAzBvt9pJOuypNjcwnzoUup/T34Ikwr6Q3K3dNlPxmLmQM4V8I4SgynWRIJfJ2Xei
KOR8W/BzeO47eSEFmLEeIC6NbMyKrtLLGxQu+5cEOXkwS2sX8plNIfWNCxyMGOfKAXMUueZuLJ38
Epjxdba/yjO1talBGFIW3fn6EJzsSWgHlWaRbzFOylcUDBGgM6GD9TrsU1R5kmBM3qX1aV/wddXk
3uJiIDaFJ04YC1FOKgCIk1zOWzXyMaH4SqoxC3EiWdAc5q3wVsaBMu1IytDYus8x/uTVjuysPgY0
ulTqB48rLumyydtEGr85q/8+GysNOwoLfLd9ejjUjbjCASUw3VhiH4lVfhi4Ha+0jfoGACLnoVMz
4JYNYqlevrX0epzsKs9UK796uwXu5Se6ZZoF1LKyOi0zcePq+in5Txvm9CD1yd7cCqdBHR/x/Rkv
p/rlSDTH9thLIRXH1CDzV241QiGroKIw269tO7hLeS7jr0J1XdALYN6/XOE1c+pRyBqHWA6sYlN6
aHIkiszFsoDd4M9bmZucw/D8C7961qaTHih9fLezZ/RZTJ81bLexkDL3QQXIBL7O3qrvTAyyJzix
M0E0RfY/JwzvDjv1jg1yny0uUOf20x7bXPGbdZR8ulLFafc3B6sD77ROz9tUDt/JsrGWjTTt9zT1
lPzuszXN3dVKOeDz0queFPAf51oHIB2aOFbSiE2/0jd2lfdH2twiD77AcPB2woSl50yo4azz1OLh
6S49hR7RdiU7b/URqg56hDkJa9sfehxly+6C7VUGpNCW63Ka0H6BGn/9Dio7S2mhQO6JkyyxbhQ8
RUp1/x5xQL+HEP5TnHCGwHgf6spyPWaz7+njMMHCfRI7KvHPzninnCIFi4Zt9dhLTvsUx5vQWgWR
NQVQbIsILVSW7AuYW8hrSZt/LzGvscMW0ovvWIwNKr8f/1dpYJik+camHZMQX4NvF9Y3l53UK4UT
LK8HZ7R7kjJjTPQdGp99ySvhIk3XSUtqop9as1FB0RxqLWpeZTSHTdOXLQYwioibyykxbEZLWY7c
TPKmjTT8fNNIdFzaMM4z39dbhU0FUgOjVh+Ow4uI4ntf2MesbAuYhfuC/J0T7l6NUQOW/VqOpLmA
GW2ATgMkderz+sp7aHPzilEW9sKOtludMGa/NEBElUC1U7j3zuO3m185uI18cNQwqoHNErYsY4SR
0XeEieJ9MWj8Tun0zMYxg7gsnm/TRdOY1d5cJ9haD1trEIvSzG3GCnRGpMJhWMTZB9zg0efuu6jZ
ipbJpFNx9DKFqHGKMfABdlaP5tHtYK9WVnzaL5p4lLeEtV6AQ4RdeDBVOioCpWTWd7DmIBJY/YzI
JSAD47+2XpO3164oUeKUEJZBPluK5OEUdeUKZ8ZBDKBUExU4BCZL1VC1j2vvLdsZxk0t2ka+MUg3
6Ssx2bXjOM3GfKpImM+o1Tz9JKNQP8jVpMJihid+7mT5CppkNUq8qbi41N5/5qYob+F9PTE85H43
mv+HWP5h4YLnAS4+vwOxiBrwbj/rDgtDPR+nIGuFAfJt7hpDaiQwr+hsPHZ2yWx/AfiWuRgbC+q7
9dUzKvSzOkQydrn9hYit7SS0XPvgZJQoH7ITFa1fkg5V3I2qZB8RCZ972IUaOoZ0cjTR/gLRUDXr
UViKeGTakudL1KZNkTKSqer00dtqKQqkwgR8FfRYSa5CE5hTlpvv3xyIn4lGAEuDeogiC/fOnb8D
oPAbcwQaLMUhC/XHfafa4XDJAEERzqIvHEO9fqZOZBYWNo3Qf3rCntBxg+t3mRL0+SBF6O5/L/nC
wonzeTV+rPfQKMX0aaxZDo04Kwx0Wzclwo0EUN7s35AVbUNqxAfB83F/6i47jWo3YswEVJxhNkcP
ykyZ4aBtqMwD1i1msby3h1T/hDnvqKaj27iQgocNLvzx71Q1mko+g8woQd5HT7T8xEjvqzzvSiKK
hMAPn+MDQ/c8SZ92bU7uReFDPV4PWLpAWKvQeTOVYkc4O6OlO+KdG2FBT9l2v4PvNrNd8CRJuV6N
ERPH4IYIcBIvjVM0yJel3XuDXiPzg+r93G6b54KgWqSZd7kOhmuBYfBGSYBG6fI3+dkREpGvUf8A
V95biz8aKBtJLmM1BFPj+20RQZaMlid3UTsvDe/ZuLL5FuhSKQ1DkY3uDDb0fJhQxUWFg670gaXn
/6tKJroWPb9nZeOcb4ZvZI6n61skUm0kCPhzU7y1P4l3tJC+ZK2SMLabJALzbHf9n8bFymzomrS/
zOTgx8QfSugKr+upwvwTqHfm9KlfvpPHUfagc6uuzUcZVn2C6pwvFrybaUAdUZuX4BCo7ItfoEmM
jlwZ5QnzC4F2vUzp6nv0P8o4NryEB5xeXcozFrmXRqZsmLtNCEupQXwIU3ZEibfhBdK8oJ1e9GI6
jO2MQKhR/AMIJji8+Em6xz8tVgGGH9GjWIC8/h3uD5uaUQFYelnYIeEUHhLrja10lqkzO9voBrIO
dNkwuCtCcjv31VUROYNTITPUuLNK7lIByxYWzMsyXd9yMSPuTemHM18Ci8tmbt7tSqy59hLViBh8
7HJi2pIxZneIpGib3nfUxCkhiKf8AchK3EtiX7FEqavzKzhq+R4MhVAB6twYmCKmgBhK0bFXqckC
SF2KT2Oqibfg+q9A47xuxLJGX0ET4OldooU9A9YRDqUcCJYAzOFU4/Dp6F4zBNa+ZLLTXbwzXEBt
18weU9++SitJ9CL3rN+y0DB7J+edPhTwcz/k5r/dtW5WbRdUQR2wbqHC3LAMaC55FEAelyvhabpY
kqu9hd4eABiMG/kM1mATCHmRoE74taaPbSFghe7+yyp8RmvvpKVSOxG/E/iMp4LLEepjx6QGuUmX
1UTK3mKXVBkVny/Tz/1cLcJSTpy4wK50ko15hnQyGOe55lODVFsB7IIOEK7v8T8fQZERq+3XTrIb
EKQx8S0F0xPW+/hIuqPgvihis9Jx2lnjhV7t7F1LTerhPPGdWJpe/hGEM/zLY4xYobSolD7I/+K/
sPXr1RqAuUCYHVWN+KJkb9iL1HUwlZlZ5xpCezxbsngZsMkEQ7mvt6/Pyr7tDqJ+y7h5oAASUWj0
MJRBuozTTkp/SdIeYyifI98iOTt83HhlNFWG8jhAR0QNJl4jYx1EIVZJRvGWXVl2Q1XXG12q0vd0
fStq1UWRuwbahuuh/AAcY8Tuz/VeoZe10NfQBosmP6wVP5y0X656GCYkwTTNHvGh5p1/644rZox2
+a6x6muInu36TyNCXk/BYNG2DSQhFJZQ7DFfWBGeiUHKekZWnAaXMbFZZF9lPXaOoecrB1PSc643
zIca7YB4VgvlznanvSUrgsKim+sMBscZy4l+szN5NaBJtoN+aQCz/ecq3hJcfinqOzKFaNv3Zeov
HI6hVXP3+OkGjX1vZMb9xuq2mhaq8FLbUoQJTxMBk2CLEqG/St6sm89AenJBHvuOLWIm/gAeBDD5
3gJDqX4XpmBgUeAkv5G2FVmtLjxI2sqzuyKK/8FiGdtNeokc5bpj84IFt4CLhGH8lyZsxc/BL4Eg
HdPGTZSWia+eKoX3y8L9JfEzouQTULL/V2Nn5VlMqOsaSdNyrh6LQXOma5j8ZhxEzOeHns95WXAh
WNjHLG8oDMsc2pe3ZvFLHlpFutkDkI92DNOBeh0dMD/ASlRoeA/E8oRANoDUgXv05yCZ+c0cReFi
6xyWIo2LhWnx3XYSEkbtP3Xf/E2q447Aaxc4pUtrBgoQep6agh81dgzVi/HQA7JtSR3baZnyALgE
BtgKLA9652mZZ9QSNlEx20R+u1AjfL9V/znBQi+zao88ROTW+eaE875fRPPYFWaj+s00Z9vvjEJe
uPqasEv+QNH1SUtOKu/bTfBWxAfY5YbUuf9dDuMdUT06Yjyen9s5M05KTrDZVhFcv1Nvdmtb8cu5
gwILjYiJqP+W24P7wPYTXwC0NSR+sGnl+ED/2Hs5wox9jCAAyaTVCYviGhJ0PkPXdqDwwOOOpfSh
6kgp6TWcSOVazJpyFt5mO3whTirXKmxi0U4VVVQ+9PHrHg9T8XyyjkYut5YgJQjFNa5fMzGyZiTj
7q55gQbSwc3jlknVsb2P5Euys6ZEkgiMmoX+bTlQB8NMTLYCGml1oN4uOGGf+Oa2t3h3o3fcgO1u
spWUfTpB1OMl+ndXFxufyw/Bn56JNDS4kpDbJ+JVVnncJNVg5o8qv0p42HA05ZuNnhlF1bnqtyeW
Ch4DzNxh8BAWZz3Vvi2FkPD5sXv/pf2yCohJTY2q2zRUZnfn83Z9rCIj0Slo+f0nM2++H2aT+tjn
jpjovKnPG+3i+XVJuhQ4BbAyqTo9xh4NtcR1D2rpEgid9KucafXp0Uk66QdjUlZb6q1oeuqVELZl
fuDFbnEThRW9nSSynztvAdIAP0YSXK1SflhYJLu3U0UpByG9118y8FYFY4zxSl9PTuLQ6tmPTP+F
jIGbHDfsXpfQ8529wVr+rNRe97TqVloNsOnjkY9azjIUCiCMjWfM3JArvoJCWOqXuXQwfrKpUQIP
MFF2aTUmutlvJtMsdBFkegFVUVIH1apwO9NrpCTHP/Cps3TEm31HactCHYKKfpvOwK4qtAFE5CMV
i5TIKo+0juNIHMkLyMALKgotcUhqpIWx4Hmq5zXrug/DEUl2/D0zMJTv32r9O9gU+bj5OEqXMn1Q
eLJwW39wieOLOB4pM42wZ/7/bkVS7b6o3ZEIOSkLjRWSi/kH/CVDQelBoz1rtrTfr7F7a4QgoMs6
k0E2u5b3ejPwl5qwkvYZuUW+FPy84yzJ5FAQ1UHmqHEV0KcJ/31NvesGGeQ6Zod4qxY6hHxCROW0
5jx+YgDZ02S+whNrcT941qYfpjHVbI8OorGhAqdOlgl/zMAjN9tZEVGC/0fe4O4zTO8hAxldDwGo
seOjcPlMtIjxNbASiSvwSFOLxgPdHecBnOngHy5C603ACQ5wu8Ii43CGVB+8eHlhp/rFtp0anqQP
yMwKj/eZrepNOigGTmvlP5biOts2G7kbGHZVdngZBDvx4nkMFpNNyaR5WNNB5jtwncl2/hjbbTNW
Ud08UsOUC/pUyJtCmNAHBRztvqB4o3Oz/L451wyZBA3eiz7IX+8TNtnY03OICgXtfXHbUO30Mlw5
fSMMXJRyFgzTqA3/B2EJlN78TYJvguuwtGBe2VA6ZZWpWDWWARShfUUGuTdC+C1CgzLBQfeJpEL9
RtcXR/3m81gxaBGaKDOnu87arI/tFNJm5dwKRlRsJXzz9xAmXGalbrB7nPLchFqyNjrEFbQ2Y7vq
Zg5qceE5SfRZKpFyJeJd9Lpke8M5AOa+ixSgmUq09rSyJlRTEifAWfnAfwIOzPzxe6IFs/FA90Tz
HM+NlWTtjcT5TOa2d7axYk5Q0/O35/3Wr3XOKumsObh1Zwy26hU3FXpeVCfpy0M1UsFO4P9olxFB
84Y732nRQ9cdr5nxpZyPNnzF0FyKIzyxHtH3294dzo5hj47P7UYD1HN0+fOWEid3t07+QFYQrCoA
xOw77HNDD05yhGCvZMUFKYRYoWmP4ZcsAYQZ04vE0M3c+fGUgpToAegrk6IrYNy8gz2aM7fv2zqj
Nrrhy3e2DZcqPAnK2DTqjZJnmt2ukZ+ny7HO1i+n29Fy3sXL7KFMVzNzKHLpaNj40eYcYFofqvM8
PM8wGo4MDTfQC1Tq5eKwyz6JjXg2ACFlX/8PcZo8C9pyyMS1ck6MeHx2gzTVjRGgd9j9Sfaf2B+V
byZmWLK+GzJlbZ/LGfwMkqtnbX9a3uPtcLtX1a0gzqErqf01senVgXxEc1wguJ5neyQwkEL4LyLU
DG15ZKanIxBlT2wDxbPSjEkAcuS9VGX6d5rGKdaCmfUKoITFcA76Cqfh5f6dyNNYRZ9aBJ804H6+
EIhAyuFwP6XBg/k+aKX8kQWX0ygRBZT7cY7dM8wl7FTCElQ1bEX5mKdNq8E394egksHm8Z1+ooVQ
hKIaCx66ztVzmMFpg6Db9dM7B6WObVEwW2oe5nKlXziuUtUNM0hw1Q/yzrKINKD/SsCFRm0T/cRc
Hch3DwemlKXti5Ugarpwe/7qq+s+DQ4R9HTbjUc8h5/6NljU3bRiKX+SfS2CtfTaZNWOkBwUeQnm
0gDhCo1U+hT4+JcZVOqMHTZQSpAAb/yllV+e+Yktnya3eI7lILntOHhKa5cGI8Yqryty/gv539zn
ATSCB+NEn2e/WKmYMXPkDZUm7/UeWO+vquY6Azi+6QfX21jVISOHVZ+XXX/Nw9TyftuzveFLOeu4
aEPC0n2XdNVSe/ecfq2mCObEIjXMurS81+Zu7NEvesh9waYg8zSh3Blt2dM+HEt7SnHFcD/Q3ztU
EwtrZHyBVG1a2csd6yY5a7hLOOGpfZd52emz9Fmt1QrQ9iyYkm0cqRxsfdtVbbi6+64GMsjepqWr
Zd887JmM5dbKtQVf1s4a25lVwSvJhcQXYP1pxSURbI35RHp+s5H4M1Rx7j8rNRGZedA15mnN9D0k
Gkh50vqUokK5eyQg46UohwgzlVOzHK0Aqxrqpn/LRNi8CJl7Gv2qMdtOSS0gLE8MgNeRhAQCgynY
YP3NsYb8Rk59wEUERorVhwsHnQV2+6OPOY6t4jLeEWXLoIvSYNxwB3mT+fdf7paotdFm78eIGgy4
ECpqr6Ed7D1gq4RX9zsS7/9yFDbhaqvzTz7tupHqojh0rFvM/mrOTBMB5hj5UgJ/dqG28TmSxTnv
HDcsa8pu+/agAwUXC4T5VMRuRyr+wu3TIrlV69G+iKN1X1bOhh5Ysdl8hToYb14sJdg9cfO9fR0g
tnqHYuSU3AbZve8In/SBP3vzGk9SsFlEXKl3mWGtGLHADEdhwV2uUNmWO1MfpEjQ8OZuSIL+MHWj
1fRM16DwxIdm5i4F+3uIEg1WJKtJd7wHRv/Fj4uC7BBerSxvCZ8KUD2P/bCZlRubDUWkCT/3gI6F
O7IQWUy7kzACSIfNdLvIcqLGf0YZov/EFWoxz4CSQT51ZgjbHZJ9pTtiHnx8PHB+bPv1xSKlvgw6
lrnS5Vs7SaNP2jYZxzqaWb/CUHVT3QOJM9p18F6oqR939uoULLitYhYrKIIGh6Sq/0VJTGinhCXy
7xm4ne5qNjSKPeUGZvlOO6QlBAXQ7bBZj3IKrapLdmFWtJk5j9qrBK2ACDJgkBVasG+268MVkA+W
omdV48EGcAfrKKwVyHgf+32F0JrCn2dFeDKMMYwqzX9jHHbNk6xCvV+CmtbpLDKOYCBLOxLrfaHC
6W3AY1jSRvOAE13tH4yOILvkZBN+qJNU8v0YcYVkifQ+KCf2dX06otiDRpEdaaKFBcdqRtBMh7oz
/k0DockUKUVnT147uHXX5UGGhhoR0VRSeL/OnVHZMraKyktyMHty5fQOkfHpYs8kiQztsex8y1U5
iOBCZUhNHP/yIHY9RgxAHClrWfCdzRKuKT3nmsVGuF++KCw8dTvLJpxXRphk889bpNsiyQZkxw6l
V663NZuwFoSD8Lv2zUmL5PaeT7yGZVnytkBhaHeBLghsr3u+sHlJE7HLuNcB7vW7sWuxQ0Co6ov2
KPKAGaGvI0BjmJkATcCZt80Y5e1XZ86ZKrhTw+cM7mpd3Dfl/xxmDDvp4zf8Q81H7GKuFFsJW0vE
odbotwQ0DO9Yojk1amqnZUCwJxRdb1WX9PHT56/x1G53Z3Z9j8Fzuf5FzqcJ/gG7VmHVClFNHOwr
e+7P8goAkvfT+nA2uv5Zl6vcAUafTF6Fw+vkGsSrITYModDtHvjHyHPBRsNPthFQnEgGfewlDICT
2w/uHGzcegi4FaQ9wfItQyXMyza0smfTDOtqGRj9LKL+w/0x415tlrKe5HsDqi32GKya8ajPcfD2
zotAIJZyaXFsipXTrrpL0BhYEX1A4ul+x96HRWUTutQigFN8nTfZRKBJ9XO0in0fapdijBT8T673
E/YIivH38drxwSysgaaJ0YQV2SN+GLU6LxFIK0ncjrb6v0mLFMwA/qZ2MXe3+Ta8I7o8AEkFeip7
BXIPl91HLWTrnDq/Jss37D5sGiUfmtlLSV331pHDbt26MYaD32yaEn3X8RWFyEmZvcoDaJmVusmp
kr5QypUqC9kv4brnpJnuUEig628x9/EM+/X764f6MoAiq1v7LsuvtwT8f6kgc+Xpfku+PWRKSHYF
pRNG7WFuon9AX2r7iSBr9G2qear6r7CDwp/kcLNlC7AFFtg/rhjxXHwrnekEOhEdTVSGOjDzO9vA
a8sy4YFG9oxUQb6lUnUhJ0SPpk23rCCyHpNGVv9ufr/UeG7T4K7VLrO6dtdzWqMvHlx1ZM9r9GPT
Oc8VvbwrzACWe6Qj8oGeN2sajuf3FXUwAEUmZPBsMdte0CvllvmBVh32xB2icOt5bK5VI5w0D4aY
SUgARh7k0IuAXcID1MzeI2WG3Dc7Pp21m9BZkwhnQZbaccbSvpGaxMnygefUypVwO0PAsOXiWDub
LpFoGwEyhC5hX2I2MMPuDnlU//3x93ABf99N7K1sHqx3f50LcZblc6d6gaQY05DLbNDZGYrP2u5B
LJkH4yOruSMYfkh3owv519bPIoVt815LRgUXtsPXNxD0rAPDLkBkFkH0ZRE7uZSRZRyhCFBFH7r8
BqYQSz9kkUDl1mBkp/liEYM479WDyGW1xeFS0f4OB1noAycdSs2R0VeYGDBYHv7zHb7pWFj8UFjI
h7Ze7cqnD7WVRG5iAbnmobq9IUPYEDIAyr+7jToSiHIw0PcWVdOLCYY7DQDBwAFbSmaWehSe/bug
ffI/nQNkB5U54B2pYkEwNiQklcnayc4Z5fXV7MThhNgjGKByCjxgJj65rc0xALZGMK+bx2Dmqhr+
Y6ue3yVwIaiQKz9QBdbSucZaSb0tuINvtyVbY383N15WY6BD4o1tL0cQDzGLfXmxeQx+Judf/F7V
jGonfs6EgOOkc4Ni/8Z/LAEYqWQZx3CydyKeR1KIwQG2zpceoZiPY1Y2CoZmzRRZtjB2mvcA4ZIe
TJsSdK8Rgqv+EYrX/Nj4q7q8Esti34eyYWcJjUktN5OzPT2ddvUdeQv3+LEnWyASAiRyCO2AJgAO
j0CZrGOqe0glLpIK0HaAp4t5cuVQfmg5oVaKLgjd1DFgGkfgbqjaMyQ3gPH2H9ea89UGAf/go125
h3MUJ6Bl0DyltunWYIdecf/4QEh9GIYJeS2yjLFBMV557WxNW0DMpWFdLqseYksFk+xWgCF/EIhg
/c0VfBvtaME5IiTaUdIdnAX32RjaH3czi8Cl9pSaP3QiVV3GDzRIkLwla/t6Wb34zSZMFcCTc4eU
YjyNRm5S1Au5wH8z7j8lkhhwJrrQx5H65jSmHZMHe+DrW2dRTBwz00uIbQj7c4ZTfdUawM0axhpg
2yhSDYTiDL9fyMctoLs09M66owZi7yKcit7eeYKxInRW51xrReNdJf6rtAkAaLF+sA+drMrBbAZv
Nk1sKq8pOb7vf0ZrtgfreB2iEoM3qi8Wx5YWYUjHA7kW96KLdFr7ajfqKPxB12lW4t1nW9JCSc0W
7Sq0zVLawLx1HdhhyieP4IyQcMhzJC9LaFWGA7yxFSbFm4922QRvq3koOfY7efoZZx/vGlRp0sO/
xKRVZ+lA1+0bmdOiIbbJxmV66ovNQsq7AquHfSw8RccUrHDPe3Vd8uwevkwX1S0sUeL1n8/ueN+8
MbqHyV2vyMvYNRw9j0aZet8TFKk4ZHHKwkT+pI2HmgmZEtFeNnHOOQAUSDyXnzAPDsYPRvM3ySg5
e849VqiKhwoOIdRMmGQ/JdE8G/JXQRcWgiEgQcxXRhyYzx3w1ISNubIln7HUj7E3VMis5Hn5UKDX
f9iJ4+sGPe4wtLlpGS9/F1OQqJ8zbVcEiqgaRxyh6X1EYmG1asOVd8wKQlTuj1tSYiwJDosESe7W
00d5vu3YSvPh8eEJ48v/ZxHKMePsz8CHLci/c3P2SFG42oc26b0K7h84aQxR0sxRxGBDLHGAN7xl
H37AEiuUrEggYC3v57h3H+bQcqIWe6SczNd1vgdw+A8BnLjr1towWR7PqT/DBRmV4y88TLEL4ieE
Fjge0DW8Ofw0JZudh9Jl5NejxupIRPdpAG7qUPlM6tOAlAyUwv8psYAU7e0GyXb9NiaVt5UqYlqz
c7EysqDZ3c39VhL20NwWJARBSbVcMBsMSYjZD0ZK0HAiglGMfTU1wEMu3cGGWatOq+F2Z9pZJ5fN
GRq2fliV0mItUtrcXMVWmHE9NxVIy10ru/J7nC54bu5DXXDc/H24Mm8aT/pTC1WyOAUqv8Ixm1SL
hlCxShFVV4L+8pPzQYetC98zXWjMwylboYmGf+Z2G+gYavVTV/7i8+FgC90ZfBJje54n/ytK7WJb
/LYcQ+MHhStQdQMZKSlgn1p6tJ/Pqs39S3/av13/MLo4sqZthisyDU+TI+YERMuE6Oqud0ogMLhh
lVKHEbWxMs6yILhHGvVH/oHaW7lcgooh0z9MZDgdZwKZanvLDGoD5ocFS5b0EZZWcxxNUtEsCSv3
10xkvDQ6Mthi++JEODp9BndRbMV+CfMJ9eNFY2/BuLBye88u9se8bFVGRLuvBpfLif9lyCGbLAOL
0viQHS1E7dyLoQK2IQVxFLWmW0e3E34m8o7Bsyzvj9EyNREY31OToKzg4s7dtlaPjEdTemEduofO
92GlHEbEcCR7QxzAYwqm1fb2Q+K/xizcVdKxWFruKx0EiACmpcGAFEBrICuO/h6oSKC92Hab0VUu
CvYQhbFLJM0wQJsCXyHfbV5XVcPDVLVUCslGaE50raZDz/6IM1obcreuwRIUs+kw3QI4Vsi8hLnJ
It3b6qNo+lgD0edsjpak7xX3nl1YeKrWWSdUwKEhvV+G3Yu6MeaQuzyRz7tjU+92xCzqxf/oh5Km
V206zO7ikG9y8XHp+XvwTCUOEg4tO9S7HQ6oq2f7/M96FHA046Syb92XeZyRbhHpkk7Wr8xhI1d5
ly5z7CrMwB8XyBn64IPcim0qmqPOOvK7sUuN1f2zVCyRNFuRSv3MVh8jHflPKVOrqYrrIw3xswab
6YFb8NR6oQ/PrRg3o1snNnvbFT0t+eVs06SZ+dAqOM0BhMDkC+vB8v8vBLRn+FXug4i8EaaNytrg
eF6obv6uBYOBaZAvBJl+jHz1XI+BXXx6n9cBWtuo6Bn4MVow2To3fkg2oKt2k20eplAVDFGYO95l
UjQZxWU9LIPYn1dDS7XryKndGWPrA3eKsofmQ9rpSgpMm35ThbLm9sHwqyfPEXDOD2aBRPgk/stI
a/tmnSqz1ZyAwBl11cxaVGJk0yVuqp3KsPq9c7a+DJOn+HUOXavvjAAVqa/ji7cWY9dBEkwzaK0I
bj+5dUpPCWwt8yyjg+YNPy1dWbeDmxNcfEoNKsQ8xsfl8WugnP9U4E1ILn0bEBWotRosG4ckG2Fa
DBmGFqPf1jwYxqpIiY/hiXETDZcJcnuSPfJQKrIYB7PmomeWtLof/kh2L8Xvh8Z4dSc0fRXMRgmv
6PjWV9d1BbPGw/XrGDy+50boRrWzZbRJwfoOBPj1IGQ8HSH+qfkEV+apdSlHqPcgaBtP0rmU5zxg
+klepaLnGejWU9CLXagjeKU5C2ek8Fn9FHge7sqWlYA4ZGxq7jzYMvQ87z8nWVwtyX2eZSbjzFmO
xWwtZz0Rt2043U8naw/+/Hdj/n1jPDbVspdXHxIpnGBfdg847sqyIaNifaOT++lU6y31kbgLnpxe
owGUvGwH6qIQVHHz3PtEA6+IAUEaGpMEJ/7tz3qT9xFSrMFN7vzkVO/RocNuSk0Xzw3IGwDFpaN9
e8pWjGY3VABpK4Kd/4vDc39KbourhBhXCPM6w24NzjjBtJ8CJIvAD0QR8Fe9R8PHCk/8TMWRHqL2
1YfTXqBz2E1UYdLwaFL9iQ8jGvcEVuG2nNqL4qqXd2SjPuR4PeEtjHvdW7KhlquN6Si4n9AE5da/
t/7owgX84QOAJ9XCMLVqo7xGKF4zdaymVgETifrtQSn6b3/XkFhHmFbrMqyaGUU7D5UUdSXEnQvV
pVWGk9R2bHgobKtuIYAhi0rkIq9ZrKXTxl8He7495RFWSGAT1uT1RTwc8Y8VIvekkRnA1bITew6Z
kvC99wYg24IMKttOv2SBadjtWIRjqRp2vBULpzsEVNI8j6bk2tPabBkVU+LaEAJBXkQj3YmcHvli
xDk279XVLL2zocS9R9ffiatYlCg+75lgv+QBVxmoPAndIYa/FcSlsDdZpI3gpFIeyidedxvGyRot
B8X9Ud/DU5j/KKAEXe72PRHt49zn+HQ6oBtU1rH3NSRY63enmlZCgClSxnyhFXUJCHS0tzaWFu99
dJO/FP/r25VcQPkUUBVokwwIw7VRWNsDR0USu26gS3vm+AfLIRMFEnZsHir2twUHL6HDzlhKP/i/
dvxC5UwGQERRepWZlrbbtRYrk2zdJStJsxVBkxHMujMm9VK5C6Ssl4q4T8kBJs/lvP+U4Bi5LNQL
SXZCZb7pd3NMjAHfvwVracMrsWgUYu6fNMbUTQMbHfDwMG9rdgI9mcKkX2kdxjqXU2G1ecW1vNsk
HoY1FzQxHzn5wupfsDHVwP0yUqgzAyXKwtKugerz+i6eZ8weEQAUC/AERHTEXi2fNlN7D+3rszUu
XCN4G1SvxslYbE16YQb5n5uKjKcsMegPcf2xPzdyUra/PuEW1mH0864yRf1DeEfK4Z4PUmTYGbtc
G1d3WjwKC0v5nf5i4x/2F8sceCt95RHD0ENHBle7bgq8pW3C3UWS/u4h1cRwqQPIa5PlteWaZY0h
BJxEMuhFP4KAe5XA9XBDnY90CYQaWE5lEIPrgHuprQmjM71P6RD1Vh+lGPR+KPsVoUI8zIlXA0nG
9qovckxwWwH7eN8zfNMQehd3F0z1+NjHxxhhDduYbHp885x5gboixchJzLcq1Jm/GQST2m52o4zq
OwG0tj50YXIwlUmIX0hhSCyV2LTVfXyZTd94IOchs2oHloHFhxZntybCfBH6/ZLXO39opYy3NmzG
JnJeTsSsE68RIN6l10HdwKOceY5GIRcCQ5hW6slZ6Qlo7ZA4HWHTKZ4hGsfK93/w+QbTxfTvj0T6
weO7hlV3//LV4VkOHpMgbQXj6qZeGA3pwH7uLJM19qOcepF0ewCpSmTMyR9MSXMSxV+wSO/V78La
XwTWoYMw2mOrYI8CUh27uiL+e7Uo2p+oyw1lcKiqXPYTC5u7z8UZKPKeXIbQjS7gp+YdQxbWOD25
xVhphHgfq60R5CTOq+ACu0eulKQvbU3E3BN0g8PbXcaH+B5Xec/mvJiEWPPqmbk3RpvpRhl63yjg
OpD1iz5kqQhj+sWFe8ahMaTCeHId4jcndI8zaqZRIEtOzj+tuKbQLIUOUssfZ8DvYsryOuVRHG5n
yFtjXMzvqn9fgi2wWifOWWipvSITOLnAs5KioSNVeYxmr9Qo3yyneCOnd2SJmSLZYP8AsHVNpZrh
0R66m7/glcieLPa8cz0ClPEVDr1JSgoMGkS/wRLqxKwyfJcSSrYptHsmNdyoBDtAEPNoYnf9DMpS
5MqN7yHwUTUdkVpxgWh9yTfk5nwmjzERtJXVOMUs7uzrtGra5tahkvDJfhiZ/5ROLxaGV0Y03OoM
tON+QmvDs+FjRftwidbA1gH353PmQ+hWGUFn1tKgcK5Zbe7E1UIbPcGGfNa2ElmGjOsg7dJeAJ6G
6oI9Yx+HG0fYAK9OC8unaHxjUPV0dOke/c0/lZsluKX4H1rHvwFvQd2V5zP2kExF2EE1QJm6uqWe
OrtKVu62vIgO9oZY807FjDEUYZV5gpFf1Ru3qSgt2mAeuC20+jZ3RreLlhN7Y2R5AGFeZ5y8x6Ln
xc3eWwb8pN8Db3VKEN4UEPxNeOX9g4AMGXDn49jZ5fUVCdd4RxOnbpijba8DAxIb7pvQQjHOwR/o
LTNwv48vfx6Dl2d5anEh3kGOxsbOKSZ0w8v7KBKpI2TqjazJ0H7DzFXsPjaQiePRXpoLUGcZn+Sl
0JFsxZj2+U2vRbaBg0eeHaI+2rKa5BFMOPIrs0b3B2ZbCXKs9ndthHOTQNUo3y6M3+PRFmK9ml26
t64yWc0DH+qlAC0tik7Ukj5MmbM2uISNZ/9RAwHA/5kEXrE9oqxwBoUmU5tjWg4N8l5xJbcdljWs
RQEoBJ1ILEmFXDtCeL0AheOPKRpjOieuUTfLzej+/Huu4hGOO1u03vI1V3mflqpHtekZ2wZphDGe
SZ4hD6vXsa/+CK9fZE901gZZppTQ5B9OYzeoV/Rmz/xevg5v/55IRO4HPFPUCSCOPaBw9Q44Y8DB
Ngz7OZ4puolErbGdPzNC0Q601n+KP+mU8fY7sE8kFWMlwwsxzY2WZjXL7yE2F2IOqoQT+qARHWsX
j18fa6CU3B4roCvteMG5vXiXVpfeFACazU2BrlGZPUsl4xjWCYz5he9l9GLaZ812yXFLeU7xIgb5
TvMMemltZIDjkdD/gBnXxX8c7jf9oPRkfPsTHpkVABxa263ADcN9/NyBl5bxglJr5j5INFhQGXnU
xiES2tuK+4Oj1HuFqRqKcPbQn0yzB6IaYKKeafDAODOOreDgAPoflWsMBAe5yJwgYebTOIoOGcR8
ad6ocZZy1ueEJ0Z98c+qSPguC9HxT014X6FVFkz+RQxrTc15RlbmNYrUR3XFjIf3lJOxmx9gWKZu
hYF6AhtIvAio5W98zYcFX8rNTIsKa9mEeJKMza+G/A4TMeQ7SG2yxLz05OSQ2sTwzVL1cT9dvjnX
PNRnuINaKp5vuiQ1ZgeDBTNKx+0of44fQo3oZwd+FJxUS+Unnt7N//FOGjSe4QhS52DZnYreF/H0
/411xmLOfl9WHcYZC5Njph4uniG9ycN93ZKXKfMjvsOV0i2lunCX4wQTt9Potgtrwpp6QlAFgIzJ
Fr92TEapvz4v432nk+gdO1RpMZicuc8qmwmgVLBBoFbHS2gbOA7JyltZ1/uH9NytCt6ludveq3zS
UYWLx31XdeBG5PAaz2GgYV1XBhrGqbj0y3tvEt+nJm9Sy8DYc12gxheN8TjJJHJoHoZE5sWp9aaW
S2RLlFbB5NhgvW+gck36mT7BtEs+GWLEs7o1BaXh63EQOAkbfTrCXlg/pVq+4s1Q/3L3ADwZQn2F
errNUwm2s0qZGuSUFbSLh9MRqbNwBwpdPuupdESXJgu8t1nrMcttC6KrnKsKfoKY2DVKkjjRydrw
m9zZzwj6jrctBSZWJGLIOahr1Z6bFavYjigySQdAp9UDlWq1vaRg+NSxLCCQLuarwlYe/Kiag3EV
73FaxkhRmiGIah+57mbzNb7lNqad+TnHTklOAe1BFJacDxNMxuAQCmNZEBQDvjs8Yh8Z+wIa4Bzp
UB46HnG3ufZHRV9wy7YyOeUN5Na827IXLgH2Ivj3ivIMkpQmaU9y+T+iQI8iEffBIS5t1dfJimzb
Y+T2TIxJK/5hmNT3XBfp4hcYztk3Ex5r0q6bZp7+ske08WXculrkqCiC9qsEaXZ2qgYQ7dUL1Z31
K+kK5LOhfp/R13L1xf3VPaFjWCHpl81OEAVR04qN/0BwR2vcrun2EpjdTQI5GWGazta2IRNiLOn7
UEBR0VyOUBO79d0sPGuHXukZTAlJaiOglWYwiZBmKU8ZD9MTehQr690dEI1rKzAk1F4IKgwpsSf+
PlCg8uNIdy9EaEq5ZqvO8r4hoLQJJmcVCneYxkfQ1pDHQxgywNLwviM03gRZqU03yULHc6KhOTkm
rs0QCXQ9DkzO5uPRXLK9FF1TQU/KZH2gMTH/ErlFYeb3UQlgB/N2/z3CnXmcmX5S7SeyVJ1Wnt9b
9t5sf8ZxSpX87CgM9FAFTKiiLVtsCUhwBwdCxjOvxwaVjgz3g7pMlq1dVkzAMVchhbDWESK56c6B
gWXmx6VHn9idO3FIRgsnCMQ4Zryy7aqaBgOLGGYLzThcT1KKPZOpCtsjH4UVHDOQ8Ixhz1/9Y5fy
LMYTvJtu7h8S7mWY45wnMqwsObB4ovDsEupsnmkFEEDtUCXurNN8QHAZh89jQVNCM5VaYS3XXIaC
scACpNKfmll/qRpD79M/4zqdw4OMLmdS6HLWprGy51EJBLMU/YpxZs+5yqI310u9qS3y3LASq8ZG
hhcluA2vaU/3R5MZb8IcL7SYCMHPnsNp4Dm39sg6M2mOiYnwX1FKPZPsgBwhnBEGYNWHiX/1jTQd
uiMBIRsh2eq/LsoHAFEfjtq95Tn2l2h2gTMV1L2ib14t7Frp3t8+UPfhgR0WTLNuyyPQB54+wpAF
PjWWxH5Yvt93hWxSwf8wjat82Hl0n9u7/fSZ39MARFCMcyMZv3aPopgbZeeABpIQdK/f9XVRPWJl
BRVyiZGMqA274WEAETffSuNl7qpJDDGCK8IOueuQeiShlmafLio1+5NPCFKmB+oSsk4WHP0tpYaZ
jRhf10P2IQa21/jGzELd+dTEDxb4ApvTfLHONJowAC7MgT2Q7nHivTnAvLQaJdYWxZWbgyXLS+X0
+EWx+RFSPdZqi2fCMJbpa+/zcvNNYcuw3ZZCn4ZGq/GV8mFP1RWIaw3oHBdeHKyR2BP6CqDK0/53
n0l5Z+7X+K8oLqLL9Zaz1iPYJiyRFbQ8kcW3BB40SMVrS89Mm6E6LLCeoXfkxnl1uPJu/4aniTb8
cniSi1h3iBihK2VU561GfCBMDQ4Z1fswbVzO09stm8WvdMgZ37LinWr7iidYXJec1jniCM1A7NSW
1WOMoBYovFbPCs5j76oFs0BPHTKp/46agFLcrbT7JGA3wskUy0+hJPAXI1Fo9aWgaXsgfOcNSyKT
VQxWmtGG/bt/rq0E5/s6Mkw1fiuuCO9n1l1QFn58ZyAJHh28WHIjIa3MFYMn913UOS8E3MCJpd/M
lDKOqpKXOTGctoYXTkdc+zn7QEqR4yI43MZ3AoCGwPOROFHk1hfq8nAIykiVauI+gUOHtgfKmC5V
nI1vxv+gzL9deVdwrVIWBu9b5JSjMvDxJliIlVPu+iIe+8eWI62Ql5YFPxHVcbh2RlLmbnnhW34w
YyXeyT7onpbMz9pGlPmNe9ZvmOHMRzmn7uG9Knt5UJe1Vnz1L6e4Lurd7j1wCB9onfZCzuSCmqhc
XkZ5JBDo1P2svH0at7GsYDjhroKWfGRZJ/4cHYdr87VH6aCBxlisDqUe7S2jxsKxgrb6ttMgPhGX
yxyjsqSkwrEBfOmbWMTW2tqiaJKPumt2k0PZb5QNrjZowbMJlL+Y+x9yXPJTwPkqolWevrrV3Rmf
rQBq2goIziDBiH+viMNTal8xmia9aDb+s9RZdkLAyYn1i0v/AVXqK/eW/dV3a1xhH4mTfpg7YkwQ
dLWhEsbD5vpqQ/VOVJN9911NvwXTlVFBMkS/QBNCZUNFaGzj5qwBIVscIBiPNOzh7o6y9TjOVn5a
t5EX5QCKvrYpPIrvBa7ZiZ0LGFKvbJX2hTygQXigbWDq8ongxzSflWsg/XtO61rZLSGOYpHhOf1p
+QSOgD+8kGeKaDa+YAalKtwEDGfMCbb2/m2BebY3sM50fqOWeiB6GNWcNwQOCHPV1PYUWmb/q/XU
Bl3x7Fy4i4hGE0uKWdiuZFT6z8JtuPU3oPyFPT5lV9CWRJXl7CKFWAGK99n+zYIj1iaRgiN28VGb
vfQW4yMJUpEF5hKNMLPkgeyY4bLR0jP4O7EgfineaoWHc17Ds4H4o69sc3k1ktETqCgluJQfHFuT
15zmwOuz9c5vhNzyy9mhFT69cbVj0P6tu8qh7ZF1xwSojcJxUwR8R3buQWuiNVmiR+j//jkYPYwU
8SXkYxSed9+98kEr16CYqpkZ+s9mkTD3sbvOdvWodeToYcithhP7RlFdFc401Ojq8fWaWS0gPNyd
1rwHLZ9g0BsdBjdny1ZZ3iElbq8QI8eVZIWjxOkVuWoTS45+qElPX7KV+QG7qm+6I6SMXCJaOer6
uKm7XBu6YqnylgE5bjd35IAINj7MWgUmZLOtBG6fX1t9IdJQ0KV8BzHjar1gtJwm8GWeQj1p7zhH
NnSk6I6Tt9yJGCqBDLl7Upz6jTw2vn7kMKShABCcTrSqanUB/isSM7r1n3TMjGjtuZ/hu8/ShyUJ
271tSATXyV6LqT4CNbNJiODWWn/k+PQUzqCGP1Ikg7Zrbfkeyba0xSPWpx9Y3As5UkwB2lyTD2DH
+4aTIt0lWVXE/wFO5BLxfxXbOrHmUxhpNIU0JtDNj2RjPb5yapVCZzX+M7XGp2mn02OHHEn1pkC/
w040n7CzY5j8qogUfLTyoT/7IgEV2hFyY2GuufCZnbRZQFfXIci6f6IsWsS1XF5jHVOBsmwkf9PT
1yA2DDVFCRZoiVHRRyG6m7EhnhGVPmr0MWiev7z7uaYjQiyWkEa9hnlTHqRoW72EOEFLuxVZcsAk
pkG51CAcmZhRIlyteo7g6eBY2qQYPAIiwZkGtk+Is8TvRVSxvBcwU+YIpriUnNRjofLUsr5sKnRU
KEYMvFKiPeQaXLnA1ElKqHzrkDIRlASsTPaVgnXiPSkNsq+w2SeBT5SsTDBFmpnRoKU09fWZvsk/
0WsMgx4xsSrcQKi+T29wQ/qQPWKiH5dJQ2w2xXYoCYkVGNkkfiKPJGU7vGADHnhJ5PCRY0szC0N3
FpdWk5J4Q0Se2Mv2KhpvO6wBNtceWJAKz9xtNnA0wTAh01cRf7VlwTokBPuc9hrsFnj3JVpBLKBb
i0hH6Puy57cyMFdZPaE+5TVwZOATJduG3UuoMt7FKnxwv/RppsKCmQpnBKl9EOPasjyRgvevl5tb
1NE9LR0Vzx6gwU7vK50Dybsxu2lkLs0HiTp0LEeDWUKpoiO/L197gJnxd4zl079OB6XXvqnhHLl8
yhQtG1ev/eF4Tp80Zl3dMJoFItkpJqAIDQ2PqmLqH76pd2Ix1EH7oAreLJHXRNkMX000P5/EjxWt
EY40nYf9Vy0oY/RZClvrYAw9ZxJGJkWdncqiw5s2yZTlsvp2SCbwp6vcFfVsjOVw593v8umdsEpe
YGJzenASaqR4XT8EMVv1EG87rDbcmgMqJGT9RCxmXD+MlNhbwgwlxcPdy0kw4tx3eUXqd+QXdL5Y
UtaOjYMh8foY+pji8gaLpF5CotZZjo+31f1WHPJKgmnBpBX5M8N6bnCtGBJfgsj7E9H6wlYtgMcW
E1Pp9Rt1xMprTWuax45Jz3DnlZZ+s9EvLe8m0kflTzsExTKgumRCxKFuxtILn1IOndJgrK0B1n91
Cd5l3awvNbvxA3docB8HiP396yHMU6eBFSevTcv8gsRbz1Uzd5CTpk5IsufRybcIuaQzRCGNG4fl
TM2QXPK7rrDXl99YBfNPJz7vmL9fhumeeyELoTfYDFI7Xg3Jtv2W4wrvaK15Z5MHKe1FGLsk7Hy+
G7cY8SmQjGG6ny2m+4FjbzEeltwScD0bDIysNz6UjkKFHhX3TqID18Co84cbi5TPP/1s/fWA8YDp
Zpcw6+s8syo+a+EXoEtf8sovxqfLNvo9A6h/Nlwu2idyjlau0t02/Sw4UhhpIMQscqQiM2KrfWQA
Wy0Ko50qbm6JPjxb5iAXV3aABJRO47WK85AGlLEdrUD9UAEsUajfZn/NIYTWYFRexoM9NrTxz/MX
Pesnk4PR78k9b0BxogDG8/PpEwT7vPi3U9dqYqqOT0Ri5sBFmXrbStLaQdsKNfyTL/rFgNFaBBC/
q1QDPyUb4aFblj7gydQz7M6up6Lqy/uB8n1qG+8t+OSpuhCOUkDZ2TB6cpiFbbLhgTEBPkUhjtpf
GukIFgsek4p+2+YGYHTm/VYfRYBe7xmBVQsTUGrZfTf+im3fN5ZrrI3sVsvTm2QvrGi3xPT2pNqT
2dCNXq0MsMynF3krHDWhRpIn1zMyYfh2vRNdbVoJw1+F+LUQFaZX1gjzD6e64d9v3r6zMkn3CxXW
fmSlqvbc/qYE8rBqylQHNg6MI6C8fgk4JZjA/a6Hmzd7YNPHEVqbo0jotky6qWPZV4lIXXDFEWuV
4j3WYcCo6Ac2XGWvr5wTfXM7ShDFT7UktTxSs9hA+XFPYxxk2GGwTj+6af763EqB+dDZYPSooumb
EZOZepng6JPOcfUp7HVEuS6ecsESnShMG6roVBUiJHa9E7tUeCIO0ZeVCyyAM4z78Jee7SCVu/16
v7RzXK0w1YPj3gLfOPAB8zS0rG5CJjHzyBbEZa/ZqOj3iU6sK7TtoO2q9btB7hwLjd77piWYu4Y4
0jnlhtSOpzICyUOKnyYurI6+RWZhwj2Jp1dR2nous39y2fMpssURNf1q0+pz8sK0NtTK2xzmTz0O
J5UdMpesbd97rgAcUPJQTztJ78X/FGDtxEa1tSfXl1LuPBz0ofupUKoOuWpX5a7m0nL8EDCRI4jp
RIuRc4ThtLH/0WPD/oJ7sxvB6RaQXCGj5tIzw9Sn6BJU/kD6+FtNqu5eM7o2OIjl+Ja3gSouB7wF
zBh810oejFAD8BVX2uabt+JxAPgQJnXU6i9lIm5MFnq1EJuaVszOgZZBJADtFpJKuTikFDeVVIHy
qkYHOVEmZIxlOItqa85XUCraMolA3cpycRhgOqG0C/A+PfxqGQvY3l28rKZAHJQ+qReJzGqZAkiJ
A8V42RR6xuAWfX+LlTkXOXS5DcovqRY/XKMuzr1nDa41dR1RdhVEfesYoPfBBtZBNX9f7HdE4adP
JwPutaz/5aB3pJxzdvUC551hMuVGn3X5MpS23+uzOBuxR5Vx0h8rhcq1aEw1Kg/IHAKNYburlqGO
EXxrH0o63nhn7o7myie2SCAUWlzCGDcyriktwFvGkD7/u395e3zlEadITrjISXIp92Y71gBlmPJ1
QWwSyy4auTVWcd+Gd7wcGc8tv27xOmVWpN/POreIy/ORsRU3gXcn2IiqOQDf+EY8O7iufrh3NaK+
UchA6wWWgXSMYo/vefXMP27bpba8lSK2NYpsAvfEs/WmXqzvIL9Ucpiwyk34nlrd+YuSMVemmuv2
pqUbN8FYZU9szUzj4xptuFcfoXRjmyYSjGylB1ZmzFCJYRSe26NRRnx5vLIUN2Oa9/FIQKFnCPPX
+hHjuO/l/7U++CXTt15ZE9J5bor2xa2jBcVbO6DLqF2NdUK7hyExKIfOTJqd5EyIo67VuGignZU7
q+96ilIzQtRwD6wuI7jlqmUWZUaZ4COIkdRBDpvl9Xjpo3WUyRHFnq9Ahr6+iHBAdT7yFN3v90Mv
ls1iQqplCpC0oJFwyoHY0lHb1KoDy4GvbGI6dW+yS2xuXh7KTomjvzU5K9o5cIZqv1oKao1S5OfL
4i/HzXs59WkSW9O0/pGSEIPMdT6NUBN3qMH6ZteZhsZwNx3TkTu8tLnp64/MS8kSfVfqTvU7E4HQ
Q+o8hd+UD62Xryxf0xD/INrFv+pc+owsODq47KSORZ5Cwsmz6pv3RojPViTjqgvfgZSwUaoiNlKN
dewlfXpvVwq1Qrgo9XTo6JVB1AAIZDP+cf/J6eMdF1jQysmjsOK56UDCJbNUNeB2wrXQ2yK+WZBA
369UMYq/4DnxXzcthvJvd3tbVijG7QVNfA4CCzScMoUwgw3UIEyVy62FN1ZPynLDdMbtRcGG3ax7
TkRV0ApPGYZ23Rg2LuhZt6UWB4r7c3S3l2LsxU6i4Mmdh2kpT63z2XPWkCk1tuKjF8XJf8RWOs1y
Nqr0ccSZk48QsXDPdk+JxzkU2q8cyHJqGeHl0B9cNHoqPABKjcdFQ36Vx1bxzWaxf3yqpwMDJM4n
nDPt1Zz3Qm7a5K6DiXP0S9qf1elCff2f/+onTAzyaxCKa8zJZjrmSVmW06eKGMhCmOtFVNJh5nZe
aVQFfhkMhvs2SDQ29VMGxrhEAKeSqjIFckl+KNDGSDvJwHgBjk9OGHNcUK+0CCiZX+wPQCqiALkL
S51ovHyOgF3hlBlOscjKZeyb6hlNvKzelAfzBbncKYXnhj0b9Z2PciB21BwfBpcP07p0PBHyRvJN
d/kMYf0HGcRMrMKh1uE7MkjiVh+x3D3ACKjOrJ3GzYe7xcHXbc0I4q+Alc4VVaALgURD83Uej4j2
S2cvKr8hnmY8RwfhNR5kCHYbYU5o6GXXuhGWsRQCD3tH58rNex2wFOhDFYcXoYTMcqOcas4bTE7d
ryk78h4c3Q5/LrvKNoIWI3P6NBxcFCjzc80AsO3rVtqobOqbs+hIb06XYloWyB3Ho1plqAPKgy6V
qudrdh7C3TXodRL2wD11XBGr5V5xFmav7946dCa+YPumUOGP4SSSpBwl0fjR4B0MhZD+Y8xaRsoR
srjoo4f4+fdKTDSMR54LbAkSHtBQW5MzmAN5nZAVLU4jG3QNc1CS0MF7J5UUzVEsrAU0h2PHsWmL
tCYQVz7NEu1mZqBui0nVkYn4ElmH+LqLOPvOZv7if3a96sW19VptjrCDUP7XfRG2wlQKcic258Sx
ur4dg9Bt/Vn39RZ0oAWkbEQsy86SV6FDd+5B4y3LYDu3DwsfW7ukl6zIsveS2I2TOsNu4Sqzifka
5gKgGsMJ2/Y7q1nj//vj0QG5rXhN+jTdomp5EW9c0/8lMcatfGb4EGjmwVuZuDY1i0pB0qRuCv8N
9Nk7SDzQrhLZDYLJ+MAE9QhuuySy8NBxcpHXMRd09Oj9WbKTRb+8pW0MSC7CdC4boMK/JNTOUtbP
B6hNZfaQKgFq8yr3En/vAWCOIoV6OYZdn6jFKV1lE1+LSkxZP0FL2dj1M0PsG51AFjrjRqVTTmUx
/6StDSR2b1WzaX86c0r0FOZbzVPb+nu+PI5lxXtSnFP7tNLFuGIWxu2wxi/juyYGlU601beq/Fz3
MelGWKFWutPlPUgL7SyVFdqMvuRxCBPcObtjNWAE6J4KN4TywRj9cPIqo04KUIN33DpEH4D41xlD
ZQu/WykpOwXsfyFVveWWilzllHQkQbEx3w4lFRTb4wVEceDr+dajfJwZDRJdAoPhxtHIsvzal2RS
/HJGb1p8NQCCLfrl4WOiYHI34g3vPPdOrdJBjgH3U4KZLReC7oNMm7zssfmR7bLr+D6T83pkqWEG
9A2ihL7mGvam8AkYJburnSGgeUIxzOW5reYrRaqeQqCpysO7nhD7p5UagJ2ycZQ2f+ZPG2K48tZU
b1w0sBAH5lbLnltX7cKTUimxRtQwelsovso4lRF4Ij4eJXkUHOYuDkPYuUsVHMwGN83C/iTRybpS
mQU8rS/u46KmFeuqCMBvBGRpdb5A765QEHpXUOnBX0UB6ZFPHs2RVAfWqmayqxZ7BxOyA9hblySr
gKGo8XLb32WjU7/8nv9mg4niAbKHso5/V6VBoYMMeJctK9P1nCu4b33VaN51Xc6ZwmfBAXzOkqSu
YIqb1BssvD/tustp4ZmPakLemEqBPqgx2+vHp4sgOpgFAo4kIM1Z/e9oecuHmAhi388ZsfAdLqXN
9UrwBzqQXnSVDeS51uSQCuOgZaeWuWEfRfNgRhGgfuE25ijMrMChYKOIxLs7aE0Qo3oEIWLROpd4
xRIzK4kqclUpfBumQkoNeQQ3zKg1bEOeuEOBmP3ra6uxE7SBi7dWSD84q7IjUZtrlcgOMn7fMUSl
qX1lwCG8hD+KGaePNHDIEp9n+hGyH4W5fHoKAcFsFPpWLg5IWXtF/j7jR2c+f7wzMzeFbb1TSlmL
mXo5pfXxjTzqBLVBJ5ZeCG775ySfjUaDc/Z4T7Gw5JmSh1XxQWP+M4+ulgAr9PFFTVNlCUpENIJ5
mJiP1Ha0IfQIjqbw2ENNIOSCFXMIx2iGdC2gecuDuxBPlAxMeUGwDiYEp5aVaPIqAg6IYmRQztwk
BAdBqT9nPA+mtkdncHVSvYVlIxx1aGQvH8UfKH8m8LXcXOV2cRDJOXNSiH/i4KtdsK4I3dbFZrLH
IlIKR/MKehYIZ7Lnz1YfpwHhCvTJBX1o3Acl8qMIJizXSOmg2JSTUkZDOv4mr86ru+OVx1PZVUQL
UhKBgAUZYPJpBh3Xaim3SnF38Kyo7G0rX/5TIywxN0AGAAa7aPVBdZZyWDAgOUpGEQBaA/Wk5ewJ
mVsStN+aumgaWsZ4pCEF2wLeEDGikFwzDGznQoq307RY4+RgpRrjHGnpfMLekbKTQ1HcHTWFxHru
pwI6ND+oqco59KsZhUIbA6K5GeAye+VBc2cVTyC9w342L4pNn2swBZquzXhnu8aoFUiLlyTM6+Wv
98ZpYoMM2ZL/Ew7fpDftL8OBwjl3QW4havtWIWQFGjP0zYIkHmRGJOZbeCq7UjAzr1zthNET91cE
A8k9isIDR5RiQQohTYs2ATA3DzyyLkIBhO6qntO4Rr6SBo1SIy1xvTvKL9O58QZ/VhB0s4wqxgrC
LXwUBUy/JFq/GdtrV+cAACLg4JFSPyJL5kCrLYUan0MLZk31Y8I6iz851qXkYOEMHWXzvcecE0Jf
s8Spg4SyA++0zRfrPUxx9O2GbKEgKx/H+HVtLV6XMMDG8fm7mi6l+/wXDgJ2wptglyheRdaqQeHy
/ATEZDt3cPTlXr4c0+2vJA5Fi/UNY+2sctzp14+MNA9KO1ZgA3OxhUpKmjGSWDZUwmhK+7EcYlem
edguJJ5/Rvs9XQ67Sc3vVUpJoUMXSLTnAqKHmzq7KAZXCjJRbFpPq/0iGZV8DmaAP/QQNX/ZPI5C
Z7qViYiN5M3v4CJ4tpqcAklgVNCUEmqr3/UsUfr0bTtunhotca1V93lGQLsSzJ39cMWe7oU+EcfQ
2Fgjxrk26KlU6uTrOrCPxF7FS40YtaFRa8TmEouEXPIc1z8WyfyBDohBQN4stf3QyN6Fdp1Jmldi
40XnDexpqNNuSVbEqzOTEaBy6T9aTXPD72DkZdFedPaTl3CyqEYRYvEypRuO41QnSdtio4wzUwLY
GYjcX4I5Lw4yAmI6fN9yQgwhkqYU/deujZlVdAZSD9q6qARRUqtq+YdN1F+TRLnh8BmGDfGw7ann
6nJ+AQBR4lkv9uYMdwYhDW5NoV6lXa2iYszMTvDzmZpeJl2W+aEGVqKgdIyfDXN/Dv6v8LPcflar
u5invU0kkbo/zvy+pf5Xa8hr6Crw8Vpm8RHf72jG6DC4YQU2OWN8YEAlGPwBuac2Gxhcifjwoj0M
JKUn9TOy+ZY6pOGlimgw5j6coN+LARXgnprQgw9gSdgrwK5j02ixcqxa+rUbNB7T5HPenhm9kwEy
HXQXsHowuvh9xXHdZcpKSaOB/w45zCmvkOMikszdys+QkxYe8k9VvlSyxGq1TnHVlSEI0QZibV4L
+3h5WVt3ljm40oQP7rS5dPJwTdXbMQVGUwdIoJXhnh7KW6o/x0K5PLCIVPi8zGX9v8oW7Pd1qAod
U/pR54PiDDcGNLIX5gaDji6FfgnH+9wLwIzBu1ybko1mTDAgZsNcl9zPqqUIdH09q+YpYSWKDPhx
2hTRG7bp6psMGe+Svocq/Ddybb9/QXAbygVHxO//4QcSrT/EygsaEqjaZExkerJuAdSTF1HXYRNH
FeDr1EThcYmB1IQZPKhT706prpnW3VNED+Ae1Zwfksa6Zm1GkkDdMeb/l47opaZGeErt0MaVyPzf
XqHwXr1L/mq5kJvtZXXchwHAKkSozKjAMRNemuVTelC9xZt31s0iUMqtEQU0UOiwg9Z/t0v3e8/R
Qov9Tq4U3ibpvPufQ8Bmv5W6yqYRsMNuSOkQeJyHNh1mp0Ld+2+xgCNl4TK2yU5P+G/lF2SQYDTZ
ww/2Cj98ljn29KGLly6JzdHFp8ZgWes593VGwj0m/6y21PUhfwzEa1vKILgYhL2zf4DPHy/x6S4P
spRnqmZHoUzyscEbcsjrcPnJYCQKM9WJg12q1LCXC0zSGM732RCLQsflokWYmsttEdEGrdLA7Zr+
YT+a2wPaY8IawtvcGXB6BGmIlT7gn43SfDctFVHkWt+KfD6QIXwI4GAg2VL98NGy5TDjPyPc2Z0d
TE4+xHrviiAFRTXUYzIocpmqb0GHVuIeq5ro/rRWU9633HU69aG5LptWSF0eSbPCwjDckrE6aqfv
HITAC+x6Jopi96Rmyg7AA+B/2PZVGXtT3QL9NBYNhXfe21bQ9z5az9wj71Ui87NvFl+w5JiZ9VxZ
8lRvhBMhaX3TrZQ4Gucn6uwaE9YbiFtetOiM4ZS4DogVta5bumaT74EZ9IiOWfenuNkK65Ba2SLP
QEzYpwWWbGNMlvuXus6Ze4FhjCd2Pe1l4nwc0dBY84j+nnTuwQLRtpKw97o3VfL8ah2BGY5oArcn
jOTbp91esfKymoLB8uD94A/lS/8tPwc46eJ4l6I3woEFulje2iHv5M7hfHBwkmrFTnvio58sALJV
M5GYiGP/JLMjjg026y0eZisCLqk0LME8SMxhcxH/nF/s7SvLyptrYIUI1YPx2fVeGgW+jAA5lcQe
0E+LFDiShUsvzVbS3IGy7a/zJH+P9Ktn+LzcQNWQOK0mveipARMOfTgYIdf5fEZh8OY1MZJm47pV
gu2t9dGSsOZz9PhOGbq/zRJGcNjqNUBqyFfM0R8pDCeyE6/+aM52orV9IhA2XrLh0KpVpIouMglw
NPdC7SazdCsYg7vxB9VN6E01x3DZrxE79/32unBQe719aHWzkX7wnmM63UPJVzlbExalyO3Id45J
s0lm/PgFM2vRtZqHn9UHo13HsNG4aX972hXJDjkbZrX0Xy04YTNCI2XOIvH65OOy4r/glQk6QVZS
1RXVZWXAiguSCHCUL1+go2XoJ8H/If64rbx2yl9lJgK55fEJiyNnzNlBhrHg+3ceScR/4uJ59df3
3JeWvuDtpuS+ypIRB/6K7fo2S4pa33GDsGcUvwTubVvEanu/zi5NMzyuG0x6Hj1FHIXkdUgpNIY5
GoCBEP1mIEUp6Xt9Pp1cp+/3KZH2fDf89dS7/TV5SABhk10znVITt5ilWBDs6sPHCr9tCm1gd6Wa
qTwbkxt15U4HuU4DirYovegnLV/MJn33ol1i1lbaSnm0z7W7DnMh4WczhfIw9ofjbz3EGCefbsy9
0arcD22cxjcMMNun+5xeViPW0rKMyQrjKvTy72vxvGVEZuB9ULOh/+BBs5XQpSMIUq45mdiLXmjZ
9SmIoCndPl6N+yFOebXDJhrlgajOJ/7BB5eIrP3brllNGEjD9sDFcuz+Qlgbr2LYWcqan6qi/vil
bbLbKfUegyM5qDzPqkHMrjTpplOrU/TZdnNceyOMEC3WIudZ/zK3sIbBrgRYrscyv9msQHNjJO3X
3E9NUxBc9Wi7gI0PKvsKiXr4gIyrt+d35STPOFfG27giqYPheptKjIibPAOshauVDZsqmj9zeNRM
/gI0vB8OCHCGyGqIjUBqcIGwmdDz3eLNlAT/bkS0Pri0Qvz/Da7EFQnGLALEdoVHJIxd1haxlqg7
x4JTbyoFIT/L/JwMH+gYjsDisUmzwFRVqnhT0vltCnJw53oJBWTWpxS6z9ALLiJRDmAzj03uE+kR
KZUt0nLNuL+ywlR7RGBp2xe9jevBYOH4Uubk4RozXq5Ey73pqWI3J0WWDszPCIYOcrhIw5XxmP3t
yBBJz8fNSZzLfWcPZJd+iliWg4qmDH4R7y0wyDZLbo6GKPhZCGKz1+SXWQyG34ZYjYABRq7NBh9T
JcznIwFvE1PTW0DytpTOWGDWUX0gQNAqwduj1HgPII4fmT1bJ6MuFN1UQsKnBY+hLx6ae+g1fLnk
PRk5fxjMoBN5PxjkVc5EdT10TXBViasLjC0ixR554qs9OaIT15hU7yPyNKVt0th4A8xsD6ImH84P
kUW9JUIU07Rasm2BfufxS9acGeZNHK6cbpQjai7o25N85zA1RYpJMgPSG3Eg5rbW/NQ9E8YHylYs
UUrhSDGvUeLfxtt899R3qSz4oeFyFQyPoFV1ljd4Txg85oR8qyWqUkyGBqL0v0VjGpPQyIWCl6mI
hO8iuE7/2XOrxmie2HSC940ahX/ccmA0QoeHyeqQLRHRW20FaUbZcSRRguTwY0TQ5eOdjRGY8TPY
veNLz/Z5dtp+AkgPIK/GpJ4qn8TYz9UYwHKXnl4pctqwrxYtXnjT9fs3yLY2BH3V7peMGOzkj0P4
nc2QoytkiWB1W1YzyxO2FlmOwZ/4vEw7Ke/RHpgRRqAYoHj+BqRH0flhWFIHU/13wRqya7cNqqUN
ZBioXnh5JllFkDLdPF7/8RK8lp6ZvP5QckiJUUx2cWQZ3J/I8F/iDETGOuroCRelIfsWz0XR5fpB
fHkAj7a1W+sRbHFqTusHH6/wq7DXaXXpW+S+axUuPfUv6BaTC3o96jC4eDHWVLNuuGMP/aRkj5rR
HyTJNMt8sBtuIQ+ilcwWipy7xUaGVGRv/YtIlrLVs6gftbWWm3O6+9UMrV4HKMf3vTcGGbCXcaCv
fURW8Zf/AQiXApAi8870DxR12w8+isDPq9FWuXrKZnOeIu+TR2EjrfiLdmUf6dUSYyqVu7w4KLvi
jYgiv0oKLwjmxpK/W6Fhe6hXW/g8/3ZLBkoSg67WL0dYq060sVgniOVOvEXbC0XgKafsF8xbWWsz
gXGaajyl4xh3ILXPECCMUBaSbOE6rbLFBeh/bmgfED6ZkTJzSzyXfF0XYGrgJ1SbXwjeVky5Nhmu
1bM5vdDuj3TGL0Y+3n7tFy8/4VFaY1a8SfAr6Burfw5U13Bd6zewxsT8IoyOFWIWDFG5FxOjwwqs
LuE+jqORZGCtdu0lanArZmdbA+623TTqCYsLlTjpewgQU6mlwLTUEckKwyVBolBv9ra+VttKWp6V
+YiwtlQ2OBzHn3ln0ZMXSs1JGGNXkO9PFoT8tF6U6H9S3xWpSOElZiq6iq6ijKbY6dGuXRTJPgGW
QZ9ujZruGhoykB3yXfimezH1DY61WgSHIGrUMxfuxorguzScZXyA2hcwvPkvu5SgPRiDXmFPyvdd
tAe26nulhtEwmhcsJsFnDfAQCx916NDnfH8nAzCRzWrTv38RIZhgrh+pBL8dw/whGl764voxjGJQ
T9zG8CAN6MdNw8UUH0rprzOmIYguxTzi8iXBHbflsCi4rFnT9Cz5MzGIrfzZ3A+rvuSBFmrsgM88
T+pSGaShjJe+i6CfpgF63i/brVUt4Fsd0bqXG+AFYEMaJzSJvTQCoWd5doZFXfm+WMh8ETvTDQdj
Li5UiGrNtxDm4Fd8uW2/I8+0vulcO971ilu4vnO3rHWNdR+kv4Eh1QaVTUdLwOBK2riT806SQQGc
h+yNAH9zjQN0asYstrswQKqbpsQ1KrsRVzjS2F+3NN3N1qTV4gHHkZDeULYcCpjn/yz2abhXJULT
ue5HQJxeh10d0fALYP2pvYEGozbe7A8xvQowTDdU3sN5I293wzxqvvA4oZ67a4D8QScOa67QA9cF
sOjr4A/F3kQ8IN749ffZSLQ2EGdkWsY/Mim4NOFf+Hso8S8LS077R6Ehnr2OVmm7BS3HpF1hvWZ8
QcfDc/vshheQr1/dnbDohz/fzi+oJxSoOr9ZkZ2AWxJSBcEGrJYl4z3V+olVfVuXr2LzHZe+8T7B
4ae1dnOBxH+Bhqo7obXdLDO7oO4i6fOM//WapXyiDtk0I2Fw6riaKa9pD52bDGzkHve53OYiHo7M
GfFni7FsOyAiGH9Wdj/+J+/whyp8zleRSJe1vT7OkoUOpx3vTmjC1fWHHzcAkCVxl/hb+YxIgMNj
4aiW48RvuzdEnTA3s6AstOniTHDyOFvV3tfc/DFogNyNSv+siHr9/S/gffMDmqAIjyfIQDfziezT
0t5N3pbXhzh+pnhCOBVDj5jG+i8hLJYUar7sRdoCk9ugIfvtsws2XV16iCWymWbAxY55HS3m53hu
vbacT3uHrgw2ttLHwco4sf4qPIT1dH4z5Bd6kRSEq3+9m2cD6EyZBG8vnOGhJ6uArXYeKT/aF0da
U8AQCIXF8pXzN6oxGfLrALFKPaTq8BI/yuoUYCouGXSJXx8uSX55ZfcAWQky4tl59nt0lnLZk+Vq
ZxqrIRwqGTdcNYXwFPqopUsXgYEkLIqBLFO6JKGwzKQhqY0IZxHNbm8d2iS2KN6U/3RD3o8gY+H4
MAmr13SlNoiu37RzsPbJCMxqzso9TaD/uQeQfRervYDky+Z0O1434tdUMAAMJegnAeYMuFssCDs7
/IAilA+7DKf5Fl03pm+f336Y6HZJB2nWMCEkFY5CtCCm0DJJUAkMYgRDm1Gsjn/RcnTAoRwSwrP+
iIifRkD1Fh5TCDnHq3Blds0EjUehpYupD3WdKQtJ0Rv0Jr6JPZKtZPkTXoxIgvODaISDKyft/wzW
RukJTHTueVkHVjr67YqDPHD0J4Eli1Ws/4hHtnYKtCaD4hkXjSK2zVVVK3HKfbxZ1hrGlt929w7s
8fbybn/3IwMzhK4CRdRBUgFA3rTkic0JP5uc5qSEmwwKkxdiXhpYwykOUO+kIMGM9Lo+oEGQ8/wh
RRj3mkCKfiE/bqjbB88XgQTFfsVxz7Q8+nI+cTWXkyPYZSaHK3vxXKBO+d2cV9lgXI6hpRVTJ5Sb
VEcbnxLqck09JTas3D/sZj5rq232FPpWKL2ZLeGK7VR5nndTVRNd27kA7Sk6ONMkFLbp2kkZmeIi
f9rKkbj/i36udBqtTw5R2N0vnQLS9c4m1zn/r8cjFQNre6CubPiry+dmA65+hbEGpX1sl1KAq7EX
Fd2E3KjoMbwadlbjuhZApv5W7SoW2PIXFUzk3bdnzf+SUIs2Tg+HVDMJ2AS5K8xFqT7f7WMDxLEj
XMoKe3wXeIkIzJlWtSrQlT96iSsezOwNXyvWqq0D5B7lmTtx3dziJxnlXek1oKWZJfbrD0xHJDEa
+NroZhx0s7ZOB1y077AG3DaHRQHNlLu/ojYS4jhHNExpPGqkggqeX2rDjrKBxy2JBuUcxa9aqgiB
suRryaHhDRfNd3hkzgNzwqYUDufbPblZslrS+fB01hGBdlHIRG5sB4kazqWfkv7pYTSHLx0QM/te
dtnJkrDxDHSsfuQHgXcQJwSDpgas24voDqwfGSJv+WmDzaJSZeS0LyFiDaVGrgm7c90bb4H35/vX
f/rOGLT/i1T9/DM+zDzRy1YofQznVsrNf10hqGCRY068fun1sslmqBmv6Ban72w+GKsuYOa53kb2
zaloWxn4bd5FcitSbAfHFAvg+K/L0c3nrFn65yXsddVp6XEizeMf1VnUJt0KLdDZUdYRSb2l3/P+
fqr54PxuGq0UxnvYDGkCv8sNf3z64ckjSrKEw7StrSwRCBGMMhIk/Gv2gzrVaeZwteZG/ysVL8kH
v/IPrK7kXvpbFtyF23EYTToHRwS4qB592cInveSnCIglO6/xzUHyYXyR2gPEJSJ7Rm4YVCJWb6VK
nd5WyWJPLeyDwVEOzOSRffQiVhtAk7RBc/u7kq8+fQgQ8gGmmas35TqcJunvlbmzyBpfz/tqhbce
1wxREX+kztw6/jGskPOVNlAwWlFWP5uBcs3x2n3wwwEH435/IdqDN44oYoTutdLHLH3hu4LkegT1
FspJ6sQsTf47FKLG1q4lgu2cBo4zR12/1EDnnri/Nh1CRAGTVpqeLkkEh65WxlXhvExirtbDQZHF
WO3It24GI7WhhCVi063DfEOHkTBOX5iK8cxIMzfHmjE93DIXdWgcuLsSdglxAFTd2NN6BBxzG+sM
3TIUsbL3P9MF+r2NOZyVZc4tYABugH0PFH+0bUi1QBIEjTYgEgchgghftNLWm5pE224wg3yCVg9A
GShWIBcjSCjv6k2WIqcjqlo4zIKYy/8lbLj8I8LCjJHwCunEgkK0noXGfKaws8NK54HrBcW3C1tO
w93PxuDOrAbVCA2FYi5a1eGFHDyISbpdCkDBDfK4A/NNTTQDZhkBqvMHrWDM3MnX+Ap7TQjtdBbN
oD0h1nFF/HT5SLmKhHUVru95mnv/F1ajbgq2Vf4PhosXL9EeoPkLNwuyUERIPGY7F24wYFFhg20i
Ixd1lwnxhs3MsLicuKCYehdOyx4zsBFSz+Aj5O+UgYegT4Oru/uW0HDWXH6JsK6wY67nM34tw7po
ycwljsnB12TUnR7zqzF0QtH/2ZAuuyPLBoXjRxed33xM11i9fznPVEpFdq20ITmCyKffzbSpbhTB
2veWlv58aYc9E7KOV6MLzBwPi3PVSqn1ZikeuGtAmz2NYkjy1+6j8LkALjp/uothQEPr/1Sz3BbS
l4dm2/YFbofyw+kCwpoHVMTxCkch2ISmjO3QofMPZDii6o/qiCkWtsZlq6aMVgIZZOjt8SfiqOd8
QH/OeLgrwAEcTL6LGv9MYAAJZW+b7t7tl8RR4gU6MWmhZ0wKZpHBIPuHh2EWrh49rPqdMOUw7q8T
exHAj/W3GvwYyqZBEpCp/MzY/NJxJwI2G6GFZzxiyFW+/gTwoMic7CjAMXe7a3WRCY6m1B+Rr0qp
MAQEcjem3iQ54MiBgRJNH2aRCWxwuUIBq2tb2uaDtAAWbyRW3OoeYRVbNTzLFzEajq++L3GvKOJg
Cvg/9RJqi+Si2Af3I1y3fy2zl8XdGVUTGdcvifpLunQjzsTm6pTJhBwe/VsisMUxYaEM6wTR200+
IfpubBp1Z7QGMn1tQ6o/j1iKVyuvGuea2JGaVPzqJhe3i0DazyuNzSFAeg1f+ywB9J95Cy2WGZc7
kFXjeeXdKz42zaLaOtLcsPYqKS1ABtMw6RdYzXGuzHLUAdl9uw9pFxyU1Js8Ae17+OEUZAHyfhzp
xdd1DKj0srZrNKg+w3iwKWwcMHchd1Fo9lAnmGbUBz3svZhArMVjgQTlRLc6UPRfWKSixC2guG9I
84sHRxCDE/8VTLh+XEheun4LVoLSB4zyBfMncoQwq7Pu7pn4lZqLhg/J3zpSi8Bmklvo5rlvG3fH
gpyvU3MM/JozMLzFQr/YHIODMxmmUl4sePS/HI4htN42mBKm2sCbCXyJLEK2xTMifO62o6NNJZ3c
y2BTz80ALWXZPguXzQkDbJaCMUH3bS+pQWm7i4HnllOEBfYbQcsUQtdsraudMOV2uUkrVKjsPLdy
hOyQwSnVI94N3WbeF8jzpQFAnMlBQQaO0FoAu9DDDUofqIXRtoM5xQNZDrOcRqiWAkaktiKaBBcQ
IV+zRshK6etV5o6fPpgwEz5DAX20yUPUvbYMXBdRyEpbmdWo+N7BxYmT/rHk61K+85SB8W/AyTz7
8OWm9AwMqWafvBOM/9Snbwce40ES31E/Op9fa1RgEXxvLEGx/bejw5IfoVaonJ7ThyhsYzqAxqX/
owZTPI/D/fRbkfVMux/ioO7SjoeboGPhiIOsLbWRP1grw/RGfjStRljrsjxAbw+C7lbyx8ka3dTp
dRaKUKGKGMegy7yPUMMxfP/dxsrRdvKkbxUekd2z/ibImTd8ydacYfkcrsqUshXycf70rkBaP1Zw
x9vDFuQdA6YSZtqHCHBvmEY2AQIqyGMjKgbU2w9TpEaKSPheOEDo65G4250iRZpnPPNcQ27eIHwP
xhNEcMPAMSgG8wQoNsywGWbDyDWNGP+AlYpWrdJU3oXZ1SDxaBvWOkiiaT/4wMHEyrIKVdREL2yA
gnUGdzv5kkGjLx/jNGchmCv1e8AyUF1SBKy5ElG5ZJKZLckNlfSSRAbblKSi4NA6k52bVjg3c7VN
7hyzY0+0ucqy7ty8hX2Li2YXHpkf2ZmIlatx7V9jMwPTJ5ccbGnpQJENZO3KeGgIOY+YhA0UVRL3
SrSibgLwFWYyBo+XDBt5hokpvi+zM0gCNv4IDhPosU7jspYMusjGw6iTWpKedMDK8jD2dgvpgHMC
kBOWNiVXkj939mX/bxvHPlpvpHRbET9G1ToPwgGePbXosCXFe6AqOcxYfxl+iSJVfpXNhGIpflKY
m2mChzbcgFRWOPueQn/y87OTJmDHpNnxg819KyULAR76ivI4uYeO3a0suVB+vKx24J7KHa+VhVRO
zlC7FGWaNMsrgT49nE5cWaEO9BGphFLAb5Di2nSsLVThbOLJ6g18/KXZHbwUGgFjuyRZFA55DXwc
AzqSa0Jd2zJbc6Ng6YVVHgm7PtaIw/ivwkKOB+5u2kwVUDcNllm7Rm69gz4NbfEdfA3uE8FIU39G
BV7t3Tqq1xt4tos1og/k9jfMexj2i3VkcBhOAB3RV4z+vYjN0UqyngGX51+/taSkgjfBVE37EHGx
H2M41TDBvlhqOR4Eb4rZ1Codw0Cy2NYI/9yyCHTbV/S6041fBVfw9751agor+q4Yi2GzSnDVqCr5
EUJ8emc//RWK11w0KFMZktVAVYls9yY1BSSudt8u7n8ScE6qup4KRD9OqDwmkQeNkSG7sIL3XVhX
P7ewTK/barga4K2DFfEo5LOL1Wf7hqqXz10L5j9eWDmdiwKaq+Hh4b34lKREZtgUA4h6iF8oR4Lt
pa/soGH8lMlQyCw+UkqBRHEL/OIp36wh2nBV+cs+pDejlJGf4YLCifVTyODNAHHhqEHMVmy0TUl9
MCMrPW2TUBd5mAUlTEK9VUYVqhVWkoqg0t04i/ppAGAPeFxL9ENYNHZlN48xt64FV5amC99Vy/OZ
OjutVJOhNQxaPTH27ajZcRkhYyJFc7yZwjlwfijC2Put15MbhR/WRyQrSLyVX2sQnboh+5ljY2ay
zg6Cgacfc/5ugYtMPIG3tGVC0qTYguvULyjnc2JW4HopQcohXaeeXZxnUdV99SgzEVBgzhfNHLqR
cBbXm2A5eilz2rVa0kW0xbNgOqVCe/ky5njxy+xSAElB5JpFLnI4zhGh+h7Xkvi629Sd9+qlRVkV
N/G3PgjMEGi6OzOu1ZXa+PBHZFXhEknMPAktYq9+uAMrzt0RjlfVXt4ldEiJUFLidJdUzqnjPxlU
j4iDjeh9kgz8okEkUt6Tmu+YSXf/xytL0ctwTS95thcidmp5OsMK7DzuzhBKf+R9J624ymwU0RWC
AriX76DHJ3/B+GCfhx41x428Kw4ILM+lO2QCcVPM/GUbtIopLWUpI2uGtAUbQnqpC+Cn0dTISYGm
pqFoOb+xt1vMQKw5OvWV59F8FD6MHwe3Z1weAmdATIrkX/0adMZf0ETZjoaePdd97ORXHMKix0yv
Mu6Wm1dP1spiFYBLYxl5ygkhkdxbGozLZpC/h2SNo5hnC81PHcn2nDqCDeH/RJrxuB7DISlVbmpJ
E5gG0q1ARDeFkB8vIWwShZyKDjLBDtwMc1gOUfkKerzi26ibFkX6n/mHJJibAj/FJ8lHW2iKpCDf
AIlHFDaadmeI76+1oe5LFysDJCP8cMoklozUUBZ9wMFhhOXxRwISos8oC6mcInRzES3YhLoM8tmU
ED8rpisL9eslwOcsQN0lEC5Im/wyOV4zl6OaUzpmMz+VxuR0EsWXFTxPaBnV25eApldNcNhzrSvg
R+j0T4h/HxIRWlbobCD705bLZjSu7j+iFsSnvDZt8afrxLSVrVbbMreWSI702yOdwvs1k8rxJdzl
2F3jOIxH1KktKNGE1Mfj+d6TH/zRhjHPZM4GKRdPN4n2Weev+BI4O513nL0ySRlDsyOCijgxZ8IF
CJr3Kpud4sJcorMyXc1dnaZomozjFFTaxfFDVOGq5P49za4Q+VxC3B0XIk8bH7mZADXS6N8uIFrG
m9Vozmeqjk5cKHTYC5bh5Ck4tyZDTxyZIFFICIlG2kYmHpVbiBJYNil7NnuZDuCra+yfKZmHN126
MciECNUKEnL3y3vVJFku5kfU1uZRbjWfv274xdNDv5TlfEG/AZwoc15RJNIMPz64XDdLBe+tBdCY
IJp76j31Nib82y7N9V5bwdtelLoglVTxRvVisyHeOXKwFlNgWfjtMCAyDKFYDcbaMYQwRFkq0NXJ
ZjoV30GFj8iDWmItGD2n1i9k6r73c/h12KHof/wBozjKX1CyduD4Nt+Et9c3wx7hMVosS/uUeaDW
4B+l5fJsbZ47HJC/dQ5tlP66uMHsC2xVyTA8w1v5JFI7GY4e9jSOTVPkevbRTQp/8uY0ueF509v7
vvxSfE81r0ZyUgxt+TMjj46BT82VRkXaZTw4C6hhDMZWC28G4FayNdhkGyuWQoDFaQCzoiT+jVMm
8/xJ97Z/FBOjWE7R4JBZPExMBfgKtb8BbEfKF5/MVtUb8UD6xR/fwxTGCDNlXkr5IwnxqtWvlRmJ
xXYlvJBBB96pMm37hkbxGExBd9rY1cY8ykzOx7f/ebAa2DLZKyuE7/tSc4qmzV4Hj3IT9mjHHZ9I
4t3/sCQIlCK0jfl+anWthN1JXQjqMuLjpSewJGIkstmlGOOiTxiM2WtuLKeMGw1HsMxtYTNleuLK
SH3srM4HJweFPWtF7xMx3IlfS1e7FMsTtOOMTDVGulJvjiAX5sNRh0NSFMMy2yRFgQKFd/T8L1Gr
a9tWWSNTOPagS3mTEbcqGrUhZ6q/Zq2ohiAsP3kmVrrUtH0ozBOyxVNDNCNTxBAKkpd6tvchqiPG
fFHaoDr5YVIHl2Ypp5NA9t6o5RhN9QFeB/eGxJAhxcIpQi9GLq2cpD2pZhWA6dFACfyDSZ5Hut/u
cSxqevvWD2ePIvG65talTqq67XB3CyOQDXjydkJqe1V5Yl2yYoqza2zem2MjCzgP9rylWF6TCwIf
vjrHeLDTLPiSBRe9is07y9FY/rUsIhaOrBjlRXeHiFiMinHP4+qWdIPOgyIGgoR7lvu7/MKXap3Z
sFUDwD5y38Slnbfo/BCgp89rwWTj94RHJcRLql+5vvWi4lgNuuXcUJM9EyvT9l4l/OSf3yaSUAcS
A6TcwceNP/Ulp+T24hZDN0w0jxGypCqnoa2b6QH2Lu7UHfdXyxQTLsSjHgmaVSsRyjM4YlDbijFE
KqCn65vaxci5HL8sLPnm6uyuwCMQ9XQ6z58TTQC1z1K7ofWvxHOXoJNEJajZCpOaUtY7AS+/tREk
g4c9CAiigQG076zRtiTuXb/PsqH6uVsxd/UNt3Q7gwbbNlp+vTWjBXAiqsdTUmsTSEB8OYAAT/Z3
GxwVO1KxG4z1rjakcO/J5Q8J3BHm0SbhmY1RSMKAQKMRNSLg2SzzdqgUYPxSctW+gykwNBkUgKek
IDgmGt6vYzJMchs262WvaKI1pYL5Qbl0Fc/52TfzwF6ymDaiftvYZbV/HJhVqQJXtxYnPTPOMtsv
6qkSXjLdazHwKmnLHIByhwKZn2UzASS+cQZjEgPZkpNXdYqp18Yx1TUXGFZy2pdD+9NFXt5kAxu0
iu0qHo7TS2KAqv8doAYZptKncO94bT5Rjr6V1ovy06vECquPM6yHRLHwo/486OvIWR1YGc6dyL1b
IGPT9mta7pVndsUmh+MlNO8DwHIhgTEP/5g6b8TOjIE3tHc+3bTl8AsUx4kdVa+ICpCDI54UycXV
TSojtSt6/HhCVgFf1+WMdEgUzEE4hXTqVH2wbfmngeYllC3yjtnVcuOQysG+Zb1EG22QEJhxGhua
r3ffItrZPlbomP31Vh18gqKoVYO+nugLftFAHycEeiTREh61PUpYbN63LDQSBNeTTCsF427cqe9I
2C7+3L64I035sOJskP1W9adVj7eeMH9KtRvTu3K0DmpFgCFCs3LdfyW/OEF1U/bBbLY65mbYnzL3
QARMThi8Mi70AmkSJDk3h3eWaasTg74ioB21dlmXP614Pvhm+HMpIt8lh1U2wq0hOMTq91Nun/hI
I8YggdKqXMr9UTuJjF9nrXWt3ACFJ4pQOR9svrvf4tKHxsY0IAGHJpelHnTRoeGKi/uc1sL6UDX1
nqukpg1/sykscIxXkS7b70NwXrOTT7n/pqLV+vlGuo89ZtVgxTydpGQlpjaAsTPjyqQxPIv7f8dK
eSaEJ1K4wE9FFsQwB8SW8dHrxwn7Kl8gA0/Zwzc22YdAaRgzU2iJbKiCwbcwtU44YPAnVm92rNtj
a6KOwJLmSZ1axXQNPft0hlaH1+m6x43QorTms2m26RjgShtSW1mQP990BgpfOdsvIT4bpqLBW6PO
NtaoWrOlg+hzy8fwqI0LBnPvOHBjCmX9aCsTxePiCUSoS6FSpr4sG+Q3etvaYiYBieVLwKmuhtLE
Yfm2ymeRMIrBw08O6xJA7iXQCZKAMfRSe9wQNGPWbU+aVjImSA3VYMli0PIZWR2RT9WgavvNVUD7
H9tP9Hx5v9yUEnKQ06KpmZefkc71uy0WtID9BTMj7EHwDqnYXGOtB/T8/bupa/5crbu8Pk5GkKla
sOGV756R/vM+fAUtrf0tn07QmnyTKC+I4jL5mpC5A4adA0a6jDdv7e/+SAy5SrMtdhh+zdrpe5+A
3MvVYMIJ+WSChkx6V/DHH4b0OCUaaRZWJ22SUAFfZAkwUeGfqJtQl8d9UkycXF409ABKn+plxqfz
pu3/i/VxbJhQdqnEHfJ3/2TvQCYDE4iGiGpCelZHuEvRn3awFAP7DA0ohbJopW/ow1p5GDDCOtEo
aTpzXL2Oo1lbNGQv1QbibQULfww5Ije7Hg+BW8YqSs5h7cJBmjQNh/AsrP4U6DUaGlVF6cA1ydAP
QPHqdAQjTmxzsCFaLQDQX2hO50UeniKX5kVBA3bd31CvTJlWR8bCmT93vpNkzwikALI71G4WMy3Y
9PZi03rZ7mctLfsJXQ017lfL+Dtg3/t6hSf6DDCb5hIHSkLDkautnM0M3IAyTPudgDqHdjNDkxm3
5NHpKSv4yFxUxsuH1pUg2S0eSh/+PZGYxE20T7YkLzOa3vL15/NM6RLxPlmryl/mrCZDhO6SK+UD
B9iqPwJ/inja8Bgip/oZddE4F7SyVXPUS52Gaxtfuqbc7X/2D3ZQ3HxRZq54hvWVWNNu6I7WubcC
pHT9HKq73j+3KXGsyvUnvlTUN7F/Lfg4EWwJTW40tSfqLkVQhbsQLrDAulVlVkHIUJF9j19tgI8O
+aVAXD7tU2srf0U6ETsB+a3iCzrnUEXp5YZAHtIyC8LBaIpEiksoaNweemARFPFDGud0JsrjfjYp
MR6fItycpzKXvnsqh1IudDXMiyxa6ShUC53OwNB92jLAD0fJvcpP4L+rFM4ZrAomTXTp9ZtRgkiG
zm6GQkZ3sOyyapS01iYHjWZvlsyZx/dh7jmXv+ImH7QQDEHxc9iqp/aRsChwH+rBhUpiYVcob/EP
AJLUakoKfT4wWdBlbWDsY1EcPoaw9sBVRKix2NQLEp8kr7h97yhDNBgxMqwnRu9Atzli+U77ZZCQ
25+8bQJrNbH75Dd6ck40Y3P81uNrjtinIRdcT/2LNtm6nLDYiPBI8DUptf7c/keyqqCcSjsC+tp9
aBeKuJgp3ue508bwOzHf3u9v935ErdOk23yb6GBQ2xmYGvRNTgfYrMqXE9/pPmLZRmH8TP+zrkAS
9qIM+z2pj7EYksl4f8KH61Yn6SMlj+K8xmcH6ZaSMK9gA0kwgkB7upawA3hl/iYka5CV8GxmBWcQ
VcHI0cGeYiasskKsV3spLilbfe+GYkM47t1mG7DDOu6nOvlnkPCatLJytQe2/J8EveL2d/M9xmJf
LZRIBOwV554FZ8Y9lMadQj9MfzlKcucJeTpfTU1v3Bc1FJTiaTss6etg/R3Fc+gx8JobjEhAGxAZ
GG0B1BKroum/g2FuDKjdnmh3vN88XiONd93XP34/7b+abFAhOV0sTz4rrY/uPhl/SUSPXo8czE0u
3VkFIChKetabdgwPaVPtGwJR6OM9dZle/hb3i7SJT7yCl+zDwRRFtHHnEhXcYYD1nzjOpdhXJtHb
xute+UueKFhqaQ881byvT/gt1fZSFMi07ihMMndeT2eu6lTO67U8ktPQedKBO3gWkN/0oDJE+aZJ
F4lRSVBU9nPXy6tqKBzcg/MY2TUIf32ChiFpbsQRj/FNjT/NtrNFMoeQtTzTmTWT+FKBO1vw5Tf1
VhUsux7Cljzk/gvqeOsc1DDGDdklXsqgytzTlLhagm+UO60XwHzNAveqCd+l0o854pXQ04Z5EVsi
oLZdAn/URwTMK3B3s1R6dil+HvHpzoFd/mww2yTR908xvh5ouadot9B+tdavYHMOmkcgg7fGOzHB
bg4eLIII7sUqRFFXeCMC6CqV/q8K08rFlP03QgNlmJ/7cebB0kJTbkMfGiiiMsrtZ6L9qn9qR7WT
jgXjuyXXI4a+Dj4J45ZyMweHSYQbWsFhNOx7MksziDAErJnqiEXoAsjCX8uJ/dx9aWHJ8fFtXcKI
M4kLWlFFaCS7A+FT6VuHj1pubFMk6/HPSQ9B76UvsDRDBAWb4y4pOoFmXWFS3w5vIw6IY738YWAv
R9FWMbQday8+yhEN3Ws+Kq0dL+JzHFloqmofPtdGSexYXj/+0KBpLauH3thy16F/xGwSKllL+uhr
J69CasNrxfe/KAmq/eIa+/O0JQ9iVCoWLNFNYxxTqDs/8Bu332VziHYlFHsswCDErxIyfsU+sHDo
EzAI9xVfZ8jSUcHiGBv7nXI0iziFn2+BX0iQrF/5EO7ZV3XypmRFx3XyLXgcDrv8anVrafVSSc3M
4laH8eWnbZdFXVYt666dbhoCfjoX8sRn5MTyTxEvm7yZvtVew0GBYAW953dnQzFxfen7UdbUi2Wn
4dq7Qd6bT2JlKZX4k9g+vMF2VWFLjLYSNocdhr8K/LivcEbPP2qnFkSD1cNgpqlrOQN48YmXdhlr
725vgC+NQdTW0AS2sQh/MjXymhtMU4RmRAzVbaVKIeNQgNawzycsiNuFdRYYi4TSGVvNvnQ4pfKl
8rpg9jGoQ8yTpLP2H7Q+g8qHX8FckvB2U4kGaYd9jy7oau2i+DXxugosTxSm2/4X2p9r5OSEKJky
v3FsUd3K+b973A3GWQhVUNDQjUg6l17wHcx7DUCF4AGEj3MDZAtNSEOmrX4roBD3fYEGnuhexhhR
NXtFUWYF8H9kb4puV6Y/785UXb5dWpkVCTJqc0wHC4d5wbuX/jVtcXiecNzI3McKvDTBD9iy+hrK
+xdFL1GC0ipZg+089NF7V2hrVuCQI3s2KNmiDV/uvGS3Othx//nhwP3oYxIxT9lERoNBS/IMrC+d
YVxL6CnwhVOw8nS5rtJbVlBehWPe5Z8SvlvoPhTdXt9Tgxmis/Nq+9MvqlbKHAVzRg4mKnqaq806
rj/3PmisX3hhZFm6nnN5TFuUw2fVkPO03dJM7yNhnlyhcXm3j7zwbBDNlGEmFpiUoq1zr6d9FWrY
9wzbo8aW0JsTAKYAqR7BD1JkSRvZBzlQbcd+CKlFsUP8ufds1Zh1Uc5/IoFuvYZhyDuQndKy5GmG
rnZyWovWnMaUMgOa/EpYNLSmDzWD3U2EkuNe25dc/CjWy/hprhAGDrQIrtTeYUKC1A1Co2qxeSJ5
m/qqoHbgwLROiEFfgZCw2CSKp1iJ+HnJw3EaZnyAuvd03Tj7Gqndzl0D2Yw5S9ICDYnmGDKATa0N
MQYg6WWcS74vfBMt+/IJBR2fPtLuIXoCetGwlVzge2xR0DH6jGvKbalMH8GDdY53E8VamWf1B6G+
eJxToCRmjfvdNThvu36PoBRixPoxVDRqYywfgz5HPf518l50tEJYbTWliUfFPJfVfnaPCXIBaGGK
ZG69+eE7VGChjc/LYRQ88PvstSzesh46K1+uVPcHIbB2vtD7j+joLrnnkcTqWPXy1rdaMbIkqarb
OgFVPHE8LxUTy6UA7WBcUNng2+JWVcqZkMhPdlxR5v13491ycnAdjGDgsk9M+gN6lejuctCHE1FW
eyi2zMAGh+I78pgD5XULsd2IKkbpzfjj2xpX0VdeSSRe8fJ8NsmTWDmDrHxEkQs9Roi8rY5pYYlh
y0cm3Ck/rOsbPtbrML1VHHbV5KqXPdM6DAreShs/IKtekIDqqtREspfoQgZ0XvSysw4Gkos5DwRd
VZbeP+2toEHu2/SPQ9S7RMIzU3BM4YUzPWN7RKwhOHg18vPg+Q8ubgx+RVpWEHM5ag5sAKfm1FUK
f1KJt7/AuNXcFdBykA3JACWbp3ur8eSAacgGoXY3I4HwbtfTAL1igsvpj8ii3OmOjdxX+nm19GF7
WKXhL+PmvtFDZqY6vh0v3diDVP2uPJItfW5YstB6IWoT3bIxlOiyKUGlDmzk+ETeZyIR/mSfIyqU
i9wCUODPL+NtQ0OkhThM8d3EMoS0BexIcLfGJOR7/ujmwUg08ao/U0OSqfDuyr6BkPz8EL6q9EZc
CbzvAw9qSWyQxPuhqjR5WlxSgs4AfPBS0SEEdUkRQNqdDIyPMZZ+KcXneAnioGPikQwXdng7gKRe
mZrztNYZNli5kDBp1c4LIV23to48av+DzMVWLJYrY6JBxx79sBjk/oFH/btJBvtvU1vfwcwvZTcJ
gRHAdT9kQkD01JW8GrPXub072MP/g5pQ9fPUMKW5ZNzAerHGYlmag2qxUBEGCDju6TwgB2+jAyXC
70I98Uhme99mG3P7zgECOEYp7wT0hz6UdhvA/T97Ua2k1/jpzDNv9UJMYKphz6Jwu5eNY6a5W9/L
uIAhbtU9f895ikHX98J7fWUC1q7ImHVD12MqpWXKn1lM1BcNhSJupNGhLWf91GLt7jwBeVizFKAs
RaJugFKP/VMJ4xduh3RX1KfcdQU0FnZUqtSsAot2i5mMz17p377Pv5zsnWSOsBMAPDiz8oxz1UP3
529hcuxwMlu4aC2PykoOmpW3PDhB6hpY5/b9pJv26RCdTwJ2yjmYi2vj3x/jfU/kUgZzfjQvzb0O
bOfSm2bLYy0rwD97bdFck4BhQg5aoMoW91YW8ebX0olxsSmVtToh5tXrhZ5+K5ozzCZEFSZ6PHFK
O1ssteU6PpsX56FHmIYXYIt/Ijv2mVM9ooLEXUjU1pCq5joXKPQpQBBdxMiZvKA2cD5ENOouejie
DcxMxlJdJxIw//N8rDmAjTc87THr/6KfP5Fgc1P0f3jkLOFdrIGqChENt+PQqWnK77IiHPalGCUQ
rr2UtsWGP6/HFPYjZtzJdFQLLj6lW6JJ6j5UMrZXqtEWcMhN/SRRLuiFmpECDRlhRSu9eN98OpWz
m+rajHtdwRIEqJfOPZBWOY12Aowy5WMFKTBc0fPCYuZ8PRZG87AmXH2veNdweKIhyK2807tyC7K1
FyT2ZOBCQNwD32RSKF3OLplAgsHEDJVNL6JTx2KY6PHYUyr8RXkxVpAV56xeoMnJ8mrdIi2AzbWR
cnzQzJxcqDCUSX7z7IODXNpA9Oo+6oTBTZlO3HQl86n8uUyegZjgHM2dPTFy4gcBQUdePhTqTULo
wrhSdjaYrjIVDGTaKACQxypyuD6TSdicPEuTtrzs/GY5IjsJNdIitG9b1ut+a22z1Nap7LbegwIQ
coSztbD4PtfXanj8OGJQsASXvgbB1HhNEEMJZdt8EoXRO1OuqK9CpUYFg8aIGqgLQsYvr3Z0aXF8
JN2XkttTNnU01QeZCitluRQpJcIRJFoONdctLBAefKSWwCdUYp98vdWg2EjsMATq2SCfJmvSq1Nv
Ytn2UnG2fGe/5DnOdfol3nu+IWy8QOG+iUTpcKaUf5OGbTxNkjqo59FDs2lsSZ01dDQUM2I+2ghV
qWvhljOfNHqS3jfrX3eB9WFeVQZL37Zdzc1gQCIKFQ7gcn/IWqzuA7548MV91SR8Fy1Kgwk1/yJG
F3jr5+Ff8pSbcAEfzyYD3xb5oW6Oh8Vsgb87q1FdtYsfFSJwCBg+xDwXjx7drnkmepD9QYMA4WBy
nBnL8FdWoq3cngQZqQg+u1/DRIWGjUqDlMx1Ci82vIqmMS9sSuZytd567VoGIYX+M9UYyiU24Wri
XAvFOG7zvOcQk6vlaj+loiub5hVUHTEA8cvAHcnL+breakf000OGAZ3HiCi0e71vJxGe0J+Afqft
ovS2/r1q3t/+fN8W05Vkw6KDQ3yyw7zpH3UHmmzut0a6PycUMw98WS/fNSPBraFuMIZ45UrZLshO
uNJbDPdoDXA/IWaf0YFZJJL8cZiwIhQXTJ4r47FHtJEhHLgzOO7RxjhjTxeELFLS/Vn7SSI7rF0s
epnMGIgPBxp72lm6pL5o18iIJNoUfzP2lILDAG/gZsb7B4y/ppRNoUI1czzggTZ91n8kt4NNOZw/
Eq/xO6hOPds6/HTGqzkbnYBH1gg/lUZZyEpoHsvRIIopNg/D9P1lzZq/ZAwVgZQ86pd9gB7YvWio
pUu9+6PFE2hVQX4Ka5qtkI6XX0/diI6id/X2oS2lx/Q39vRItskaOF9lMPzIKvRjsUOVM0q80oZU
2CdGwJVOIQ+Eq8QGDEoGqmYG+A2TFAgSEEXJ0Wc+ekM5SjymIHGjOmGW1mEXW3IK4re8jBlm3GDr
1J1OdMphp4DygGC466txSAaz93Kgaa8QHUUdRDmvH6IKqAVaoZ+TSvk7VXbyYgnJBXoV3aYvTQea
9Lc21L+FlVq5EeYSpZr8tD5bLXbmqtXxQvBD4JJj1uonScQ3GQgwOeLuTbvi9FwGK+BoLlMt/q17
qnX/DD46Fu2SlLKk5GatGu3fpByMx04SrtpLgpUQFO1DZpjInWftWSaBgzRZIAyr9R2XmssXMnpA
AJi/HFC4Qj4j/QH/mzmx2/5z9g/a5FaHrDN+A/8WwyBgOi07v40Rr5Y+CT6tBUQ9C6jfK8f1WlRt
nrhXOW8UmFKhBNCUmdS6VBEqXd8ohfg0SeC38i5BqL7m/vSK9p0QVzMCI5Kk07r8i69Ut4QHlbDn
26m9uAayn7L0j9SOULULkZZxlZkqeUWx87XrB6ij/97TUAApm2ehPQWtGqY03XdW3BtnueD30NMF
wHbECA/PLjycmX0V4LNFreFeEqWYsWYiGcJuHpm9U0i3wKN0GZyvOzKwtFNx/wDnagL/MeNBzjvN
zMtRcvTfF3bRu8YY3QgE30B91+gCjIwQfnYlUv0SkoAex3yY0UoydMOHLREokB6Yhvz6OvmiuKp7
WV2Cd45knrPG76qncsYAkQ6CtxxvlnDf7CkbyW0IRSX5XrTzgjlxv/xQvVhT/g7K7sa9AcdSP4xj
Bebicr59sirfiyVGkNJVk5l9u/Xi1/4UVVTfRzd305ygMBvoUfaHRPqbhZA3H6NEbN7od46XGQG/
xaw/K61Z6urVoCEFuXOG5VmsBXdv8XgeqYmqyvX9tAcXCM0WHCfBe05CoZb7l27lj4SGZzSc/6vE
Hu6Th2I7lt17pJAgirQUqaKkkhBIrZrhasO2gVVBvs4jn24tJa+rwiWSA+Ctm0L1HEBwSGPeEkyR
ijvQ0H5wASOW7NJHE8TwmijwqnMofqD6H42VX4qHEA7AV7/5kCB5V+CEDmzx2n/S6aJ2gHCaY9qT
1EWAlA0HBUYfDy0K80R/49J1k78b4pGRbUT7yyjZjUgHRZ0sP3X74jODo0I1UJvW5HDVVpaUn22U
uEYI3fDSJrtzfW1SVERgxMsSeH+ttqH7D2LvXVSgQa0HZlDz35yaQZ4SjapQl1aEXMozwR2P5BWH
RCGZKbWUs4Ik6ooFh1dH5EUuWANBEjVXP2vEehYwH6+TBqsSheMpd1rhp4hb//dncgf8qRD5quuR
QVVnb1887GRjc0lsRrZwZc2DgmnM6Gk3KvYM9ovEPse4OPFJGTz5/GSJtEnpA6ODGI7O3JhG9xQi
coYRZP58blMCcVMHIRYSYxx9kEIOmZ8lGSJAWtTzgoMo/zdyom6o3sqKDpH9Fx3nXan0GvsSZACH
Q8aIf81GhWH1quRhkl/4hhMPQlpxCfd+7lCsfU/fygPFTYh6g9gHUr64ABjs9dlxVfnYVgzS/Zqs
D8aPBkTu1iBFY7tbOwSlneCiYK/sdokzg1QcfPP5mkbe+gxXE1orqMRiVOGl7o730MFpM0rjSzG+
KBoEILUEbvC+UMQvW3lVtnbN74nNJtgCOZBjjX86WaCr/2NASNaaqzT8l6QCELrPumdZSLzsa3nl
/0PNHFsne4AGZp6d4iSNHTx6W127gVod8tOT8JlpE3GR6RsHOvlq4A33ZNaf+6GxacJm6jSdnQap
YxdYRXCckJD2Jq7d8X+yKdam9tiqDMIOkwHKsPG2+ciusEie/G9Am6Cu4ET95AG6rMazziSt8vLU
K2ljIW2sBOZsEoqi6sz86flGidAOMZ1IDLCwX4s9V6MoHmvaodLnxbM2eBvLaBcAzttd4CKNBIvi
+I029Lym+NtiZ5HYAiDaH6shy04dmzBDhaMYxFz4WpfRRylZV6bcdCAVV7gW5w5npjzqbX1lijM9
hJOR7AvqHkZRHwRaVWMR/8gaZDylrDgaqHCFHBPryGR/0WAdcO1S7PiBggyg1tgUQmi+nGjlKjwm
FxuABgwXZkf0gWGaxINXR+A+5yzTPt4j2Zu7D3nQEztuziAE/jha5fgOmcXPZvwOO5lctWKkC7Eh
82wmkjKmi0m+DzN5u5raVIN/OmJ6lwp9XGYC5e3yuCHV3WFSlzUr8uocd5ERLEygpTHBnGp0omsf
duHbVm9FhockiraZ/rFiP52I1LNPUeuOprC04+1GgxN3+zVsH1C7hEpwPkl/cshjBalYmaRSzhOQ
ypH5EgzOaPbic7Fug/4IIIF4FWDjyuB1hIIme/Jb3c/ZN7i8cp1AUQRTytLsp8M2iCpLgEhoal3H
R9NR6fxnU6KFBVHbcb+JLciYMZdtfXrh3Z86Vkq0Cj0MTiQtMsuHaJcmSBynOPz/w+XMIe5hij5K
iTO/ilhxhhGT0oAu03w7P/lwp9vBH7HVJpedNZK9YNqjXvVYplft8RVpjOVwKluewkbsewXF/mZ1
4ILzu/vdFXQfqxzG1B1F3pHHl9C+kaNMy3g6UVzjB02qNBRT6Sh1QJjb/7vniAtkWeKW0hkwXKhQ
V9/FaOKCwgPPNKE8Xy7Zw1fx9fXkHfdzevcOj7DwJzbsKJDwZ7OOjqdvPWF5aXvzeoaylXN49uPx
EVdv/Li80btgxHEYFBemLx97ybVjZyxueL5+g6ayJ4kJJL1urqX3brxHDhgDJSzbIlsX8LNA0m5j
+KdVwcjQpYhlqKHniaiJ4Vnc21sYm2swcH3rjOY8tlr2eeDDpiSTS+PLltNpISVZ8gesRPZXMhD9
vU5ZNNZ93xsoWmoD1rDM0uUWRw2zvOz0d3mA98OAkUwlIBM1d576RxV7zEDKAltw+3lK8Qcg7DVv
D8p2v1C9NiiaG1HeihYkKqzkpc/+3djSQpRkMISXZ4oaoPUdcjKd3Tys+W6foBa/87xoGJMgtPGt
sp/KgP80kLAfZG00zkgG/5P+eCZv9LBEj6tlxydEeOIrsMozc2zppzbrm85Pu/KGzWT1itGo4jzS
sTCQ8K0f1YAZPhUfDGSpzop0iDlCnBtYT46kF2/0Eu4MGd7v3oo27TUa4fyLg1aa3ae1DSJ/vNSE
wFGU8Hh4pgMQOIRhD9fkKt4hskH3xKrCflv46yG7kwaMjWyl96jNxHw0utHozK6O028YiYYsiQAk
9h6wtYsbdilT3Ou+RRP+5F4n8+fcQkBpITnEezBpP27E37oe96OXYZKPVwtHeKrV4epSMbfrWNcH
Na6lxWEZ3fhPxgUIPUdEejnhnEE4kXReSHlfULs6J8wONQLG1jHW9dAW4xmcLBoPZsj0wwKuaO3m
es4SYzSbG54JW/N/zgmOseaJ/YrhgWK/E87I9Rl8dDz7LRYtnTkU18Q48ol5qYlD0tqb5qylNmb6
e4a7DEa30vinvQ3sYkTeomY8XdHrknY3niolsifmCEzBdi+RxOneQ5YEIlOZBh3viPCWXGsjEpkx
6D2o7oWNwixhK1T6qr8Vp7mLC2LNrnvsrS5CbDC6X1lfJ/p/Joabdt9G1Wno/ZGpt9JXfI0cV2Dx
dbCUwlkBoJroamm5B5yY3hBaUH6FOPQ7JKgFZEMs3L10y+Zqssr3aWRWwWQI0FCMEKEKDNZU0rzh
m+Pz1asrvp+2VuvNqPCXoKrHzUkDRwp1dl6TLDHmm9tdZxku55ZGiyWQBfsz+nI6trAbGMrB8kgk
Y8uqgT/sQga2XmIq6+BMotCNUibSlKvglvbdaF0r8eYLsE9NTmOYCeyk0sloWZf8tBKBQoEV/0xp
b97Dc2bmuQ0NA/QSPwqGn1flYZRss3fQjB9HSnietxNnyTid+XENSjCeLn/9pLgKbpdB/wDnuDYi
VETZ9SN++LDxKTwTH47gj1/E0/q4crdSKlCnraSs5dNo21CuvW+BorqiWPHu82OLfB7QaZHWHgFH
fecdu6hJ+JOl85Zt5c6V+RNv8h1MGnieaDtnH5BZQZGwrcz7EgHzowMlXulgVr2CjpXGCmkyqbXu
VBRsWBs+FuzSBcMrErpK0Z1AnVIZIRHgGi6rFK/y5MhKOYobYvOQy3FBVJXuwmhWEjhcs8s6MYv8
95RTYR9fFvZN8oFESZbRg03WiHALPB7lVCehn8SJZm+lVd6iUDMQK1u6rJwjFoz2WiUK1ToFHFDY
GlKZ/CtIrKnJoheLaZxbDmkKkGPNpi+ywR9bwGa6yCZq2AYzkSeRt/9L/p7BTtXNjzr8XUEUDrh4
FVaGT5hzsWZ4YWJkaiuMgH5FBxP2hEvmImmHY+zlwiazcHpWNw39O2s/I4NFvOHifoZiVWZ6av6b
1pZH2c/3auCBWLQjwD0n9bi6d4OfjazeIyKbV8dX2IWwJklS5LjN+s7+tvP0Am7OjyOrlTI+YJBk
4uxL9n/yssddVpWfKJhoSuP7abV+E3hf/bvkzhsC5ZqQcj05O7EIiVFbTKYLcbxrAaBvY6flGhhY
k+QnWLtNLiThQp9WzVDn0TyQ8hJvEBMb/XAN13Z3m3jaByR5kS/HcMm/0QRL50faw1SMlkc0DLOv
+D+GEPr836MeZOtyXNgZq8mIXr4rR2lOx3SAno914OjokvteL9INLI8+vFmho/ImRRuyZTdg3DK2
aOzaPYKlVwVrRztDyMgFJA1QaRL8VVcfcfvVut/1XJEnaOyvuAKdijj9bew8cDRuDw4vdGn4nG8n
pUMvj8C7IlLTQNrKOQOsfFytSn2yUkE2lSJ1uiCBrJf8wf/UjnohVaDlon1Niy1nTrSjFgtX3naf
R7LMI441AXDOwlFACgi7pZYZyUiXFS0Qd+qsSYFlHkZAKw8nytW/5+95aMF7DqPovYDoQAXZ+/3P
jjW/x6QZWYUU0jTIHiFECvxVDvGxwY329HxDqEDEuBbhYwP/3JhLAObwuooJPTod4ayTcGFAFQ53
o7I/bbDq1EgFFRF99slpSOm3Ifw2RW7a6Xb1Uk0qQsJmXRGa5YHC2Ch2zNn0aejO7S+zEoGXiY2K
DUBnVBlIQ+J5d9NfoD09633fKm0zwuB8wuOwyw8lpaiGSOxPNEjlOVGmossquZGn4ZbIbuy3OZX0
6FfBgoT81kbDo8WgGI6RAcEHvG/3K+W1XUuzehD/Lmfdi74IYL7q0d1Bs5dcfe6VTAfFqJIk+Y8H
kujzq6rOEF+Vw9FLywO+a0E9s3tJi/eM6GZqheYHnsh9W6r7P/A5RvISouXyvwlkog45A58p70vs
pdaXo4bGW5SzS2vw72F+uqwZpeyAB2DHE4A+GtDKmfcsamv/lg7vbZjzblw0QcDus5PPjL536HD0
4RaaAAYv6z7pf/ijAuWmlVwEfFq8+OZ70uWQqN4I7/7jw5WQ7mhHSAVqGylpZ+S3hIB3V8ZDB9fk
ac+1ND9XTCwwTRW6+nl+b8VTSWMxt8nQX/D2T24F6lgC53Fmm6zneoR5kiyJCLlWF/hmGOb8haX7
voS3pcQUO5V9QJHPf654yuSrfiEdZMHLNG1zeMF6Dh15NgjQNcsF0vR+kX0wf2Bh8k5u6RjDtIPy
kvwC1aWIcvjKxqBRsfFmP5AhfxQc5qt5ZFj5Yv7APrqVYbzwLUfUPmV5uMMzMxXBnMvqqRKCfsTg
AYUd0bzB8fa2XJa2ZfZjl1J9WTGsyQAv5RfrBsXFXwQ7Ch7AejPNzUFR3KrwdHq/AcsrZNo+ThR4
s2R5Qh/EnqWOPVdH+m5mpvlT9unhS772TaWs0gTWHoGpCf04Ik4VgePUyoxHg0hw+JZm+z/SFw+T
wKjYDGbegginCVxijQ/Mm1AR8ujTmTxOboMOFVOG/gK9kkIHqfs0ziGv37oPQhgP8t7D5RpnqWML
CmzHDlv/HuQ9GY4CX5ScC1kC++kGXMG4RLQMh/dTs3i8ILVKV+hMkeIcVTQlgRB/IoHcR5IVEIlw
wO/llKOgITLkFExs+Q9NgXRbnbUkMZ87YTAv7vKjm/Wze26JhyjqTI7Pl8Xv8UGyI7i7WSgdAul1
QR63u3+xgpP4dpYikYrRxZWlOC1a0JeQa6gU81KBElaxCaVOHjKz85/X8QXnCDzPC4Hmod/2P52g
Vwbu+T8eP0rGUHtxFzwPCJkfbZG0KRKsjkg1EIxOb2pvYqPe9dKAr/4Xz4nMpyIWrn8+wYQ3sSgR
zKgmyMGnFUsFNq3xNyGMnINrnM7AtjHqdSoxFazvjZBaRdlaUi68evm/Ht+d6PufRctTN37Tm7N+
MfDv3CobKPlhrWCJGVQccd+9pBewFptoFOeTJ/KeCwM3gFqUp0yrWi6Rp2p00Aykbt/hefErjr2j
EMfis9q7xHLLpHHXfuXCysSj9oKuFDKkMW3bCTLEgjFByBmLKrbS104l9ge/EDitfrwOf/luX//V
yC7XJ9OiA2oLtW6oPeyZaEMPIrWv1gDPzE2Ef76/reUc1hKKfabD3w7Rh8okJoHpKRLiR/chHDvd
itTg8rYGEGqyd4asngW/258cgtXq5LpuFZlFjyrs03F0R+CmnYU20IyCvjy3zI7Fvam2dYwDDEgU
1mYTgASXe922ptdz8bCOINMGZJKKSvoQWhVbpaJzOHuptW8NjQS9ZEp5WEbkqnJSwoEIoIFBgT7n
afgOH1meFuBKiH6QzpdRLFBo9qbb1B3HryF3xsRCOQBZEGv+deZNBLOUBZJ47ngOLmSCRKHdABfU
rHrbydv1RiPLueP2YbICBi/gjHHCVgO5y5OEvD+LpE+OqIt4oSAx4T2KgjCixpihaYE7/ArUNiTO
++3U6DFeDRERhK/23kDQSezxbVpvLiJO7Qydy3LPtoI9qn92v5XS6q99J3QsOj7Mnkk0k4epMmRQ
nzaU3cCjITHb04DQE+Kwgs0EP7YicGgp9UStwALpD7ENrquZxP7wlJuS2Ujp6Xb3CQ9qi/NWUDDT
FisZxnVpQ9ylG8S5dXbXB9RxQ+IMBkTjUVbazzK9gnZRmyBnabIVElpPKK3tr69/ZURCIXOTA/Tc
XemDcNj9ws6KbF1cBxq8fUJxFWG+X2N3og/KdyA5WkweAvPSyl6YSQzzttLj4niekGgFYGpw0DR6
QsyHCYgm7pR5ABW/2/nM0/HTmkJJt+eT9+u1sG1VvPkALO5yzQVCD9HiQqO8XMnI3eGa6eI5QSCO
m2tcOvKL+M/CIKORN83DBFPW6XWHddwb6vlG3dNfG66YdH2HEMiHiHQ+f7ojThULq/a96kqDQT8X
TKP8WRf7LmhJwFZLRGu/O3CIoEBjFkegs3jXIUNOARD0t5NG4EgYGepSfqrhmTE7Xbe5Runr2J3y
y0swaAJincWR9UVRrZK+rDfaWbgOITprdt666UkuuRQRy7E/vJSmqKQtvs/L86CgN3LxlNUJdNNE
wENvE2006l60Ir/8uWTQ7O8ddMwWL9SKgt6SDx0CcUo1Ia615cbEURkg04mkQVlbBdQ4DWVW24Xk
f22Rlt/2TsF5gWf0IU79BKvLdc79xBa+zZH7eBcQZIzrBq1m3CWzbzFT00Elp90rHGA30RfCL975
CsGcWDhgAdfwx3N21xmy3/QZ271bMNxIdi9stJvv1+jS8cURA0msYbtqSqggPuKE80RTI9CEDNPv
6gk7uJl24kLgk4cHaiNB68BSwTaMxwnI2VChNl/B97XE7UZmkmhysziTgCXrL8H1mNILR/uY9QDC
/gkKVnvTwPlC7DQ2WNqE0I4ki+oSwqIXKwEuaFjHW7X+QXRETM1tbr2fcQa4LsJdTkQffS63b8Bh
BtqyzPqWpomWjJZYAsz8jA1pUBqIcmRJDFdwz1iudwBfqeEoLXZvnIlCibrQkGGJUOxpgpnVQiYp
75zdQb3rtPMLWB0NTdax4SR9DAlZC0AiAJ5qLHN3RHBeBsDNM9HBRZ8GYc6G5E35dEucYnRNSCjJ
y66iIOM7IumcplnBJ/beJjCZp+XEk4qYEqez42gzBIC35rHRCq95zwXmymZV2Rh7bhj2pIi/WO7Y
f+dGh5AaADpZxhsgTp4rWthLA6OmW0GYIUqt6okMLvAxlxRtFjXCVOmdKPLn+XgPMMuRhYkhX6sM
XptjjQILjr4LTfd0exGCHQ7sQ9URnfp1mFYfM6no/dYBksiPuxlW7Zz+Z6RxcjewkqEwRwZTGfFl
/Lg12oF0nWc74FBkBGBwZzrJY3OW5Xr8kVsrXqpCWcoUq0l2KRGH92UcK15ViQWuW8hhhNoGW/kf
3CsBHdVeNH3kY06IzgTgqS0GcOkg65jfraWA7wnegJ/HJfcMO02mdUriHvVZuRlBA85msCptIeR2
9gcoPP467YLfUFv0iA4lZre4ufASxaw3Is5nf89KxniFo6/uU9ihRGkGGPy6PP9hhYUa9F/yfGvg
0dKhINROFVsQBLxJidtWccDDvAcPzZKO+1c1PAiSqfbmH54Uc4gSpRWDj1XD0cIBASPp/ULD8zwg
yt7jKet+pK6VCN59O13spgcUel5s4xTMc+lHF6/KmaavRNegpujVsleiE9tNq+wQ4yT+dnbxH9WG
UfK0HWjybJfr6xJmWnxFXNheWzDh94B8A9Gh1KCzX7KYKqmewc1cYDwTFYZqVNfEdW+Sgh6jeUDl
Pd1aJG3UK0AAhirzFesCnfNyhA5w6x5Iu82AcuH9CEU3rA4KhxxHQLY3+2jDIrGtWtPAKmqHKKdS
t1A8ZnGrNw8dBieVihFUFxnZQR4sp2dCrMoVDxZjbhrgQj72Y20i9Hj0kC34uA2gdRX3y4ZWLtMI
ydZK/odEbEyYhnEo9RlmtD1mnP6uMepGtFxmyJceZwW1MWP26MfzthbpdwYYRyh4jtabnKhQAMUb
SxzSuc62UmqlmUbU9D2xYFuY5wnCs8ozXiDYQ8fSFA4WiCqFH1C7HT6sqZBp4XeGc0pZrHPy1+Hh
pJpcsumooaticWzBoik9bIeLaHixWMZVXjpWZkLQ7h5WAzYdtb34Vl24Nr0GYaTu7J00jFUfDrI4
zLByJVSxY+8TuV0IWJtUrVIdPkHTaG1lrpc66RbhT/rfVxNSSgx87dg+eTm1PaBYk1QmrYD0irmV
dMsYWKob0BqJeJ2cNFZNL+lS4LNO4dMGVHeT2b3Nk1hBPkk6G2IRnn1B3Pn090XJQlU3toFl/7eG
YTOi7r+0mB9TD/Td9O2gwhSIsBWOmZUwmgXCTe9p8DB5zpwF/wiC+Lt8LLs1bJi5hAR/O3THXzls
Jb31l4dBbveFvnXivpH43dT8bJD9t1pAupi4OMHd1jGzVV2SINP6bQZ9unQFMywJPE4aQ31hcZQr
SxZIIpNVFpW37E+34ODL+vwwxgPGZ2VNYywlcxJNFY0U4RoWnfKw4x6DDlRN1NcNaL7yzCaJiThw
y0ds1tLgBnctEcDgLfzzX41dIdzoWnyuA/p4MM49DG4yph3jUNstATqijBwdURvrxlNutgVI0q6N
aCaLYhcNUYckgnsgqqxqgoZNmHD1ucpj6L2JhyPfbepIBcybCRBLmKA729ptjN9STBIZriGfHgrU
+Lufwjv0CzTEGfcGNscwBjChP8lEVwxzdT5XX6f/arTtBScO1jLexqtxzUw7kQ5QgB7LsQB08l1X
/+uO9psCuv9b7hogOKaGX/CLmO6Ia9n3Rv1EwvQwSRemfMTXRlyPAfvc6TisVmQkW3xqIbqpb0Lm
CyT71LahX4xC5qiJ07U5Vb1tYzq5atrW8nJ164wjK1abb07FcsyqxgrZ0SnTGD6XziMgiwSovvHd
bqwtakhbTGk+AZDL+bpUsmrxsjzjrDEz7T4ZSpIbJprpI7pTFvwGpYCOeL2vLJyvsImWEM0w8Z1Z
qs+f0S8fIMC6oW0W7RPs/Bkpmx9dozW7/yBPydcbEo+X3G0IjJHl4UTz5JjAmTtVuOgxNHq6sNnh
7C46MNVDUcE4VzuiQuFw20T17A5ZovM8ifVACwqzMHFmWNltakbU6xpL7WVnpUqepbl1YpLDMt5d
BNhrMv0n7KYdPb9TT/BziTiajK0ronK7C1+GxIQpiRKu5pKs30AIYEDlN1JEhKRKTcsdQGbs9M2k
VHGtcX1n0k1+XcwO9knoV5JdOjWot8iOguwatCuc9avkVQMm+7XoqBIhqWLKXrUwmSzT1FVS+Kt2
dgxK60GpCn+VYvq5csZzeeBsrVHgENuuo5evx7/N4ZbXu47+bRgQDnlUCVbWAnb8QryNU1ypAKsV
elmwIz+g864bvSNeCLb3eDmvJc0O8LtFJreocuOXdmzTDM37PJYGidxG9IcjyQZwMup7bnBdacVQ
4mVj3NdhCmt5pKIPfcpj9rMZgV/EVJk8D7ZaU9h6ATMWLalPgSjwaJwvCa7OUSlH7EBiaIM4zXQU
OuGxps32rLtdnSZhmxJU68pNw5RluLdsHRwbHJn9w/Fm0ZGyIi930O9IRu0zEX7S8hReq93/eXQI
1x4fpRyHM/+bSJ+HgB/8YwpSZgthuyUE/nYru+sL0zV+MIxwrg7frwKoTVMDwv0trRVXnRtGxuUN
aeeji6kSAlXPnEIZBdgTfxqPeP/Sz4nzig+FDvZfixIIMuBab+k2uc9aQ8Ux9u2CLXmcfqeRwIo8
9c4OvG33vaBZxJNAxZw755PI5PrX4Zc9vZhuk8MSYw8tRPTZApzKFo/jTOO95VX+oVjmqAV7annp
tA0N0p021FXdwfDV/rF5UavtM/EgJHDO9l61R0YyFACbhFeLdVtlPC2Bvr9YYsH1CFsJpsxKR++G
Jl6EjVC2+TsvTNs88NhQKR11ZF5fIQC4/ENYdm8YObM7964Qa/NeB+ke1VMKLOzWm4lE1NPMiNH4
EQ+ooCPwQe+5kt7Ch+42GRzP7sMuJSu3RNyAJeWz9W+xJ+obVnGjDQfb5Qr9mmxI75J+cCXSmu2c
k2o+gy13ZqRoa0An18elvItg42TLWvroTr0+PDndMBn2BvFTbHel5nLXulhp0oBaa8BUeL1xGjnm
muhI5pOuabbA5EQbIYS8h0dFwChcuCckpdEdWs0STwPFYm5hoTS7uaAtzTBrHV3IUS596fddMl0D
jmAu1F1+rsCsRiWTOVgVsHOruBqQ9tY01C2rJPjqWkQbXJwkobfP0ZmGvZXXmepl6pF3kuPVpBRC
Ml5mKnoaR/sg0XKJvhq8PdO6KPMmE103J99ZE/vTeI8sBg9nmVyyxs47/8yuqpC5Fm6aXYXF/YGr
XRUYzNzj0X2ERo5QhYuj6+1golDqaGZ733iBbAjY8qKQPmsDUZSlYdOE+5Vf3sagajyJwGzoatHX
5Wv9/2oOhDCjVV2oAb/wq9/vjaRM2+DqWCueLvS/6aOROrHHLKM/VN1QCGHqzrdKUgbQ0WKmxGBy
avhAItV6ivjvyhGMszXs0mh3ebsf6aU7pIQP0hcUS60X+sA7wveGaE0fbtuig9FJpeQsTgs4omU8
SerWoEo+xSrwL2PCKFxT6B8GOohNtiqtTO+dbYmoBR8Pq0VD29aYvRigOgaElZmOykn9bk3zLSTU
5WGp4CZ5bXFtKkQq5beSSGNIfSoLnu9JPGmI3alv7JRUffOIvblFGmfPqdN64moEBz3vVd1875ez
ecejc+EUZeZNI3+mvi8oOM3ZYJZTI69tCpuBor2Zd2mMTEal9Gfia6Lwc/oN5+lbl9FaknD13BGN
0o6b+Ha2X7hwar5llPeeEU7zBS9toMOrgA6ME3QkPs12+khPwoS6/E8JGPFQw631FVToN5AWXjzp
Vlv1doMjkD5VQlJeuBpIlmvTEk8Q/R7LU+hwP5I6YsLmZOIg1Sx9rmGQ3jL4CZDwjViHL3uJfB7s
yExAff515kCRTHOB/p0QMY/J0GXJqMu0dFBvgsrge6VEUzgD2OwxpnjuboMt7hxslCVtjI5E9Y6F
ehRYTC+MSVHi0aP9yctqkFqkXD6ynfKDA7QukDG2317A68+5cJYo2TjarbBlqdOGQB1zSThmj7tz
wLrUjWfTkied8rsu9C5u8JxYIGZWENILDHPLkJroh9cYSZ7XAKKYp2+5WXCztVrOGHzNitZq/NO7
BcI+3mZ8SoStkQHe4wolFTZGd8rVUBt0EsEJS1zhDWJAIbdZZcVCThuLwQGfB2SgGBEq4mCf/bZQ
BVovc6k82bUtU/1r8jYv4+eNEagUP+H9iYyCTmP9RWxb7SIzkuLCpb5LvhVBlQ2gPj7ibk0UqHAj
8xYiRMuNSTXYOvm4hDl2vqFsAAq7tfYJUrW6sF0pKOsw3yYQObspPJqF7o4Gu+Yo+KT4JrN0IeZV
bRNbMc+/WVVqT06IgvhyKlBpyf/oN2kluydtcM/d3Hlq5lySY2N/EpHJr4EaO6Ij7ftCiCSHI3Sa
d5JJBrbH0nSm1Rjluv1LOwPft5Aiq+RyivGA+4wND7DHvkUw8wfD5PwyWqVq6Q+wo5zoBuicK7Tk
aP6rvRrHtDpRnykFzcRolIgmFjzMfYZR98YQcv6sB0670yAYOT6c0uPndiyCUwBkjlspOZE3bIBq
4bSt/+XfpPB+p8wRzO2Q1OC8jf0Kot9GI3ftqIN9FndNLnh3o3IlwCDLHgoeXsy61CaCDo8sPfKU
5PYE52dIRllgNEqCIU1nPPJdfvz+banA2VMmZ6rV0yxXPEN97erYIydFDlche5O/5edE0ujuCYv5
cUmLJPCeVarQgggLoklwkbC5gkw08UCyGUjpkh1YZft3m1op3JIjf10YomKOD3awNCPRfv7kzBYk
XVEzkYdYbqVNyfDKsHSNhFfeUT+D6IFo1vkX8EvIq45eIrAfh9pEueMcAhNSulDJqDSEjqGLhK/W
O+7w2XxKvdrqN2rhG7BU/w2+rjbUfNinUbF91DvD5doTma3S9ek/CDMEzkCRjb8wqAftELVx1SPa
zEisq1BUMmJK8NYZ4ZouheYINbZOkWG2IkNnwAWIB+bpqb4v2GOph7rGs3yzQtfU62zX9ogvj2Af
dn2aSnnhjKH8fwVKtlLRqPmGDO5L2vroJuZwBJ5scq4Xd/72PSqPun3SGQHXBLCKik6Q0b/TYufL
Tn+7jptHn0JzATDehqad+uy4l2vynjiUpxdCLq2NFtZ1hswS77uDt1cumIF0/BCgP6CG/wuYcnix
et25mu+7mudOdbW9hsVQTlECqixKPdXVe8pX4G051zYPb76ld81DOPdRTNa5zADCdcAhXxUskZLj
xEjDknNsROUt9FIcVIqlCDZ/8bAXVwLSHJRiTlIRjqSY+L/MJN2q5/uXblmfEqDl0rqyOyWszuiV
806w/5ag4scLmKYMfYq+tjAac12unDKWWiwOn3YGhGB5xe2SuwgZmnriiFLYTbpbFFIx0Ik3DG57
WS2R+j5KaAEfL3muo4vHBBnrcOfARSY5HyArY00HplQcwZ0cfVHriv3uK8qomJmLnbRa/jdsord6
m/gh1S42xSp7jpAjR41AgZ8NHUvQGy8u0d3Lr3e54CLqh+yh+1W01sweB3dOuWr6b5vV9U/kFNOW
4oeOKGJBp6Z/4Ec+wls1zyYQhYZs7jBU9jSgYsnoCiAy8pQUf0BYuGuYDjywPJzbeB1ZjZ0U4Szr
gZVh5ta2ANjzgNrRBrk7XGEF3qU9Lh/PUQW00eP0hHj+1tAdTzp6p6sAxWKuEzbAq8RPrvO2uM1p
FByXlbpf33ZlKvqQs7Eqjw/Rg7aLsRBeEIbuwTIQpZTpCf9AiNISH8pFlifa+vCZr0bfGl6y5jmP
D1jHDT7nbjDGBUqcSdQj/2sTcdHQu3qUu++u5J+xA5O8f7W9tgfmNSKOuQWWqrVDVu0B6wHxapLV
NL/gdUWFIRZCT46gKHyBVf9/uSkoUFeGjt7ALEHllo0z9+sQLfbBxvTqI+SpS0ad64z8C4Ecqag9
Y7FoDlFIbtB5gJEwWvgm2gAxzAu0TC2EclDlPaa2tfjd5KUqzaY7L3dRIE8sPGqPt/X8MExCl2P+
qCEjMsTIL09sNc1h4ccWRkzvNq0GcVKyNF7GxOP8JeHn0PKfZXcHtRhLORhegZl6egG7ClenYyYX
wd4vNsG91aFCf84QEaPTzuLdXEy5ftkW2tSvb4fGqxmPWNpBqftf91J59aIsdWm1EcOVFR+U9hjb
5whAWcuKtCqH9zkabJtUY3ox614/IEU8B6+b6TyDlSR1ji7UUuOEbhryJ2t/+Qi3vYDKvM7qOmJn
u5nN5wkdCiUH0Deaz+6pPFtqgIBfv4AheNgfyCPPNlTvAxUMZEvarY+VoCcIfdwpsUnDPEvIYDzm
+PiM4jyaEaIbmnc+sttAEXcAlUhwe4x1ho6FPrC+fTyYvG5NPa4aM/3UxWym7597EjKX6+KQgt3z
8gzRcrD931o5ijwFokKmCT68ciMuk5Ub6yAxg/EwcV9tkPobwDfGXGkxPbNyl1AqgXFn7ObTfxNT
7lQ5xG7MXXDWO6MF9cy3fO+jUdAezQN2+6Su0k4ZeETOcuTEUkO7F8nu2yTqwYs6OMS4bQk1BHsz
Rx5UZe7hVRYY8iKfAWhrkQvexdXc948p7NvGWc85+d9dH6JBdZTcDtWPu+2ykZPHeVnXgYOOiNTC
OmOhjZdTKG+1oYagZJKlJ60PFZ4XYYxNX1YSmt6O32gXTywradcNdekh3BaoE7QaJd03TPcRASnq
K7hmms73hiSCoB9UoQtmfAulbovtkitOx9mZGazciVuWo5hX++dTCEj76swullzANazuSPI1v7L8
g9UGZpXCQUYxjksKDAd9Ir0P9heefPJFBSFhaT+s0uufgg74iQRM+hXgcdjdH7GFKz5Zu8dy4RFF
oM/wgIb0BxAwOpb08IfPU+GergpQ7DR3en4rwwJ6DPDm8K5Ew0viEXf6Be5HwqhCGKlByK/Df3Bb
SPongOBL7Lm7ysaH68UDt8sDhgzTO0CUgEksLms9h4QdKZprybUtCY7dJvE1oo6vCVJPqt8CPGl4
f66pasg0Xg3wknAS9jzCsSbMmMz6rgzGprUk9FP5W7ngizC+k/AWzQZaQKDLys3mmnwFznPKumPp
Ug0eLOnhXOSWSZqT9Q+7HRrWIVzt/pHC1MoR2T8OeB3XAZzylRXXfXcJdReumuOkJweuxg+OpAa/
qG+7AdaLOe7+D4AFZ5wOWhn8Ce42z1TfnokwkdeoZfSHgale/EZbCQsOhoVSygtGgWmPNYUk14YG
1LjmOpXMdjerR6ZXgTxDcYO2UdkVWF7fBYa3/eSyACdXgLg5YeaigU+pUBXe8Jvvbif+Vy16x/i0
yuz5fy9qgxLG/yqTsaUd9QsoWNRTdrK3J3DEUGV85RJekCUKLaHRpA96Cmdhmv+2KZXoXBPxO/qi
SvCJ0TbU+4ERQ0rvcf48eM8lUzzGGSWhRcP5ijUpf7ot9nbJp3gkIvpv0FAWs95DqpCziUuSiZxm
Od2GLun0Qi4nlrWNoXSclxUxjpvKBG6XbGb/a+/I4hcj05YgPwPJ/g0U5ktBRnNG9kbFg1dZF1P1
O6DAnewv7hSv48/kqluqQi+dBugK2m3lZmwyuPcMy2libvS72sTn2Ch3e+rh+ze+SMLrqZSMQLKl
sAnFK/H9C8CmENZ3Qbc5tPD/cRxSBqHPhWbtkcL0M3Jv+67HcLKmm5HBP1dzYqcVb9ZXQpC2eWto
3Om/wnNYKBlDT35+GFrCYigOjSG6iaLGFQ/RZ7VwJuH2nNGWldcnq+yUKeH4xRL0vt0pGvniEP8G
S4AgMyGf28NkXCm/qNveLpfpQZnMlLYMgh/iuADmvYqpCDYczRAiOERZsK9vL396S5AmFBhPCrEz
IMJW+VnBoSDgfy0w/OJ+25gGEwRt7HAsKsJ5jzEEI+zzdrtdhcI8HH8GQPAnOhuFdoDvBtwwi932
OFC+8OHHmd1UMlGJGwnc4Qqhr8t/QSre1RiUAjr7ye2C+lUTy2kg2FZR6LV16DVtAWDVm/hXS2U6
b1Ec5fA0cbveKdlmc2Gex7uGukYCXqyIu5f2FANu2X5GtOR5nm+D9XrfGgrW81JCAzTSUzLGWzcU
gi+wdyvvGWQasuRpL3aiaaZv88tHUgOfVRpcEfBA2xvcLMQLGpsCJXtRw6num5oKYA/JzrFv7Idz
joNR9jEp38ZxM3+TDh+EUqQIQMX3LzIJhvRmwD4ru5uOd1lrOn4oeNq/htQXxHm5qJFZc7IuvVS0
2r0pppXulsqdjzf3QJa0dQiapSF6MjnyPWZces4Q4bAmDLNyAVosqjs+Nan9+tn6OY71R9Q+Ful2
Gxrdpsf/iJwIXw83k8dsBFuPfpxrXFfC3AMITopfoajD409MTxfEXqkVKPt1iWqduehus4e/47BN
lcJmBeTXBOSeSiwb6b84qcwlasBQWPB71PlDY+xh92I8NlTAPrLcMfIQaWIa5z1ocCAZ2T2L5dGh
HdNltUnDRRoGaTZILx75j1yWSqNwMG9DkWe7IkWB8JPZsDNOC4Z3FqyECpwyhS29/q8AUiLafP2X
ssNt2kAJYbB4C2xDaZNXKhj1ph0aWQCBSRHwuX+RTVQ070U2/hc7odaBEfvUxiFiWx9Vv6lR6UVB
vP0J3Eiafhvpso24kltH48WC3IQpV9VCFc93updMWFzG7+VBlC6y415EviIzFWnAucUL4z9GszLS
cRBjIobsUp3KOrtJGUmfaGQr/O6XVJ/ol7V53MddV7y7x1LXZTpSkLbUjl5mNEflsyguKfnr1pr8
zdlwremusVt7pCq2f2xSG5q3p3a598wmHPy51HN/6hcJVkwjH7yZ/frA3JkT6dwFq+jPuUMxg8S/
UVVMJXOtYP/Q3dueScCyy1tOE9KmZmUzPcezj8kfmvb0oOvHDhZAYn3ZifwtX7/VWcdGWNEPotQ7
B3PUcTawKMf16sMYRWvx/A4brSZ4nqfTdtdHg5qllMnew0gK9LxDj+jl7c3OxdSu0hYO+Xkf1KV9
MDlP3FaGSp4wvrtp+6mNPPxLsKGnVBojj9t6XBNUOgOUNkqbAlbqFK2Py1wgx8id4m6kUMJGqffG
LkhlC9FmZL5ICbJnYXlNHlYjlauugloR5QMupHitAX9pfR4lPoF71S3wTK2rtJvkgLL3QdMNlSAD
f358kWBTAkwznyIbCVqhrXKyphjl5OZW0geCc9LGkmlgJGcf7zdUUYfpI/6Z5+9xi/a6hZoijOva
VfUfOLewcS1lDhl8nSXpA5jdH+XHIdjkul5s5qO3F+KB2Sf0t5OXe8mSFckEhGZse7uXXx7HUIy8
3wWeet0Yrk5BFK6KiEsmWaTWljheq9bkd1siTpCp/UcD4ELEPc8nS/gaGkh3M54UAdiH4vNDrqKO
yAlW7BLKPiWCpbyobLwLwbjaIZgowx836Ob0acXFRJ3tP9ZSHmtLm4YNcw+kxYtJuoDPy1Vo0TFZ
XNEAaoR7a7gmiVlzAwkmxblsV6hkFBeiRMjtkl7j5m2v43oNZS0PTSdLZGjUthSkq2I90sjajB4D
eR59SOsdeUfsSSW7FYmZI52w1hD83YTbuG2iRCsWjUbxBGkzGC+8AUpdSOK9hlBtxi3PsaS7hElA
tEJxEymPQCMNn9fvkKqPFFxFebd/fyKoKeI3ptrWKdLv47a6tbvKfPaDa0ejuakd7NVsVMCz/xuB
LJl1tttXChGebk5TqwwNSqmbm5feo1EoD/Ewnx8WHe6O4ngAzvhunnLZof7VqzcT/xTKCD9LJrrj
Rdkuvk9PXeq0AfRW1uU+GtFfVN6HlNvLWyzmW3AFz7TTDhidhx7z9ZNOnmBapSGKgFB4RXVNnxTD
xhgMHpJjMyH0NE5pTjerXoFUl1mUAP0CI+YI/l+HfEYcbvZ5MEJsd7Icbc0H7VwnGsAeYlK+d7y6
g0Ssfndgb8CclnfZMbP45OCmo3hBjBQKKyoOF4Jbxp+sxpRgYXP/CUWMXXVcvGXMPJW35zfQJ0wY
s0Y97bg1L356tanNThP57nUEpegOxhbo94HkK8MFk71UpEruCWjDXZcnQfPndlGyCs2OerUW1Iv4
gGAIKbez7SYno8P5csmFSaYhSiuGLSzEunpJc/aAo4DpW1r2kzHxtKLQyoTJyOUOLnGRShuHiZ7G
AMUjb7PuFKXBvZ6r9i6BJyK5nTQF0HKUPrj1vDSv4erlRJv3DVOYrLG1KaugIhWakv6tLM9vMeWk
ffWYQCQmQ3r+9E/5ylQ9I1e7XhQRUIC7PYfsuh3Pz3+HHyBJ2CPSZn6CcBpMtoCPewZU9FvVy8A2
m5TxxEFJDChDLSCELBkIcYGephxIrYEXIJDLIcXGo4rWglwJKDK/0LNZQxS6TSdB8rioanO1WO/t
gRqvD5zChDjYyQnJhQ5rLRbd2LhHXLs7ZOnGvouAUZRDdfSE8POamm2/TMdAMfknaYl9KdA3MrST
VaMescg2GKgmim2AjsJcobOYlsq7s5s3myflLwfSrNFdqzQFRD14kq7qaFPhAfYdxI3Wx71u6AYR
QHZEsf20NUNK2IeS4U5DT0KHWq0qr+SCHWAKLLi8ZPDh9U37VQjkWxDCMsM/YIsvJyq8OZw0Uw59
09HriSC5PnIJC7QmHdrUJE+H8WLzzjiBkpwhmhw34ayC6rwukn/UTdRA7Gj36sd6IMG8xkUtkjZg
RhjH3Na3Hlk7W9SbKUUAC85uoyG6PN0C3zp35QAIq01BSsr4dyDsuauIAHqtEnR95cM7GuOExBz2
rleJ3MCQVq6ZW11opLfUVKz/yhU6ZtbEBQTOIqN16EG7ODh6Z2OKJ/llVsWNemUc7joG1szU5hrl
SQqvgMCmcz4l/SilX165BBlkKNOXlRySX/IWDsL2+uXV0zuNeL1pC2hPqkUN1nLi7iBFUDkgkb2r
riveXtiiHrtXEQ2LxPimvgn+LC3Zp5Hp2hWgQJC5thdiX7YZx6Iwun0/mBuboceVGFRko3dVBRrY
wvwjTAHOu+NiurH68yv8nT45HDJg4BOgNpdXGyOHpDFoluFqtI3lPqIMOWlnU1sZ83u36S3v8xhf
xdeFAbpEqQnExGro97TA8tuvHNIfSYts2tV9lXZ+Zq100IB+Bi+0SmcJkL57Uewj+OtuOrWkhDHt
Wb9bTsWxJgni42UBq/7J0cRFabofqOtBAL+wc1spALDrhnXSOwDuz5lHWZG8D9zJqH7Or4PdPNit
mhfys1m+F+zzSAmHEVQdB9ZU4Nh8+QfK9m7BlGMnv04ZbOnZEjVzBUZzCbBAYG73HQPUOX/uwT1x
OEH3UOWVbnqvjZZ/gjzXD744xBEybzBucGOZqkJ5/FFeO+6upWFx4SwVq8r+8SmpA2xJ5QZar/It
XkB4dlgr34I81c+JXLSFt6OVjCBPfccYG0D0ZYreOxoyKLDy0RSDkkDqn5KT8R6aHrBA+r0nrspt
+o39De5nalbA/UZr2g7Xqj7otI1dTdaE5Rvz3eBtkHA8q2EZbasRgQD00sWU1NIzaAva7Wvs6pfc
XIW55VbDLHLFS6/waQdEfy+A1iRLc8hMg71Yl1XU5nJJguWqXYCxV0ebqWQWaSAF4PpHx2Q4kvyc
E++fRehSKSGflSrrep3Hj36C3VZLuGs1IdlYqPadzaOQ4HeEbrw9vHXCCd+274VL2S9TUegEJloY
N/d/q9Lbd/1z05tsoU2/eKUF7NT3m4+3lzO4aEYKVOpId5y1aJmPOlfUUHcpNn2bUKt2Dyq55ZH+
EL6AoG6GU3rNEZunxQVbY0excdv9OmwW2KCNk7Tv8Rn3jmtN3YffbQJLLax1sATIlSVcfHZx+x4v
2KuuNo+9cDk2O9EX+raKyKiLElPYcMDTK1trC/o/hgt1QuJAGhrpVIitiFz0JLXg3PeCXL+m/Vdz
reA2qU+CRx+hgXlPM3vleJ6pU+2URjBRNuQ1kYEsWK+aUIYCpX2G9Jbm6KI5/TFFchQb6JxNjgg2
ZpTsKMTVl8+B154srWwIUFRg0mCHsRyW2uYxp8uNf9tlQ6fLXxtrlPeMpPke5hW1e7WXTE3K1E5o
Hkv3XlNQJAasRh8610tfCYWaYzbkxOJRbmcuQzfPCJhTKSaPkiCc6rW73iwGGKFpeu1MYYTBp7Sr
mAKvgaZjDsZn9SnVn3Qq9EKuUUqRNadbGXfUBgAsU3AZkE3ao7+hyvzILfhcOogVMC93NttCV+9u
BqfBcBLifN9uARQ8D0tl3vHt0l2kbGXAcMwqjO5sso/Pcui9p2vW8FFvJRRmBlvH3khc20/lBg3h
QR2qrT2Kk2sJ3BvSL7v/+PtSvHBMDfSo83eK8PRF/RWMrKZIO0q/sQGCkY529V39afq4Rvn2GUXl
HLJkfDzS9EVSqzwxib0o7AsNE44THfACJzp+8OhSkCfw/q3mi22zIdxrg4udCHwm4L57lh4t3Gii
EhIJYqni9lcTXIm95m8wBdWB6ddGkmALasVMUAx8MIdMei7eEfBTNHM+R3s9LoMA68LTbwRdUrhw
JCBaKqQcIhe/JUzuqqJCoNTdYWehG4WYcQ0JLY3O37A3b3JcomPiMefrvsP3mhAE9bSlDzp/s8Df
gjDD6XDOFsXY0NiwzejF1iaoXUxeL4NbHHq5j8V5LgfsUt3FIgApf5FgE3T8qr+H+mTkLuPV0j3e
mn01M77etIoJ5t1yAVrKtqVZcpwYxS9gsMKHRRdH2Y9m/9axy50hUIpgmomc6q4KWQje0aCDqYz9
JNQefsGs6UY3iwqAqSRGey2ZmFgdruFodWPGNeR4xOuEKLwPBsJKgxaFUk7ZWYYavwFEOIhpDQoq
MkKuomiIhPFodj5nuClT8rkj9DUZg0348cr5TMdg4OynkXTOph7L2EcojPUmQx4iDKTW+Yox7ElY
yuzBkgCxbPsK9Z7dT287oXJlDY188xslEdV3/+isk22qdPzN/kue5r4n6bkqJ6KyhNN+n/iBZKGe
QjXeb0R64swzoYVTgG8Hy1R7lqjUrA3wiy128B5457ZRfMBmAI7vUejKsQAraDoFd63qD2zo2hE3
QwQHIuJojymsHTOT11shyaIt+IQSfHQm7YCVJf7+aOx1HwlemEfJUEBTBKgf+ng/ZWgqdFLVOYmP
nnjAUGem3K9anhIgHMJ6SHld84TdY1L6T3S+1BC5umBOqE2YSMMkJtepuzDy8uzwjwZBUcoyWnFp
7OOUnn+36lNiPrg95TpLedAIyTXYWe4b0m0Xk5f9NSen1akOMlHYtMtoturdK5JPlkS10l/YTwId
XIspx987Zp76nMxsP5VM8OX3hwTeJfoPSDvBx+oF/TlPZ8OPdSLnFo4mpu9j9Wvn7AfdoDcOqNOt
boy8xNQxvL9LDS9GUvEsIZ1Yz/8sKR0Y4txufr4QMlfkZliqI/rLk+1BtrYs9iZhJeWyCSsJtzac
PvF1M84txF7XoNwcmu6tBQP720hrStUlUnFhBQfa3o+/sLmoirPY3d8AtafK82jnaBX954uRK7C7
/08rPPupD10fmfk7Oh3Uwx3Ad0kij0T8+y6EiYbiY9qAO1LnCothOTqcnaw5WwR9fBs4HUQNaPBH
Dr87LuAt3cIJlR9cha2GE9N1F67wzY8iebm4ofnjEQ0Yao07hAXEyG+q+XrnZinCsZ8E/7FtfNrN
qERLPX3y5yXWyRqaHsqt6HmvWtGsI9XZeC4xjf1R+JGllpAURsmweSFzsuy3grPv41u5Tj9v1Byn
8RDxOBh78WhFT91TcQykNja6ajResOvXuRE1O14g9AavNyZEUIv8izGWFDUpF9u/TwLSLdeJw67T
rXrFWsv2L4FcO2+fck3tll7s76GCcgkifO/d7nt+P+u4ucHVmVowOYB+pT9tae9JSZoajD0vcVkZ
yOnrY4JR2YneRcuUvfkwLQRhESGFunqJZO8sxyKCWXsa2X1PQr4A5lxS00XcL9K6RyTK/owghsHA
irTi8vUNnruBOBHcHOm8bO+Re+7bGDJNxctwqVb1Jv/BnuGtRwnqPPghQgwvd0Z+K8q0fcwxOhZ3
kcRdovFIJiQU7EWhFzCgVPgE8SuvtA6WTRpyPFOL9XuAVQYGLaBMEOU1vFrBbH3OaX/WaA1z67mu
2arMkLKzmJS7chbo/6aXNuFoVa8AtgPQTt6codRb2xSzq9n72KxF4g2j182VV+Hb/c2dsay2Q66W
8gKzGBwGMdTNiGVrkqkFc9r5bbxPqE8/Z48IHgXdz96Q8Ntcw7siYkC9iDWbcKY1UGpzvscgF/vt
dKHzdkBtik0MRixOAxSBTPaHBovHlc0lGy1FPglet86w91GiS8XT1MB+ICRAxcxu5p/n+dsvutOs
XqeVBeJlRsBB88r/EVpVxH9EjVuBYeMBRPazio4TqUb9eErt/ZW4SS+TixXcAOgVHn1OmxYPv0sP
8UNqTqO3GIvCd5XanIajkiCULqnxeF+mNiz1YztjNXa6N/czbd0E0uMRtrJ89ShUKvMgz2fnuVjn
2zRNduDVW8SFzYTYbwTkYe7QcrEcFU+YFksZdW3XFn9/g2wipjVrxtPG0y/ezeZ5EHNvR4ITFk75
LKZ7tIyT8aIJ1sZ5TUwEHXwdJL00La50+D1Xtw0bLimNE7KM2mtiJayc2y5KVU3uWf3+66wOB4ai
ATcV9VGdEGveooM/ngz97LAu3dhj19G9QZKsOXcPu9kOeu6lp1unha5MuKcFIpQZ0qJjQjuwxrh7
u3d4237q21OVA9etM8gyz5V4PxQb1lotJ/QbZFrzcYUmprpdAkKuoqKimJkIfI7V3dFA0JUcmHhG
DHGbS7b2kAQ+0B2Huaxs6fbExJNMcBphPNKNSsWfLhECRSRKMTTTVOjl9slNrj2gC77TUmKh53PT
YJIi9IcJgU33udQrIGSFuZXxxehioF8j/qETZDDgnlk6iXzRiCKktCKfJe8AS+1mAgxFCITlFKLI
QxpBipa/9G59jFY6M8OQCGkcd0ok16ppYCs3VPFvc0JcL2HEf39L8DsGG63doasHXd+p1PNKRnbw
d4nWRgiWguc8daXUa5+LZLoLAKmabzJgCFnYnWbzIhTjT7bae786lNYWb6eavHPTZlzjE/hbmzft
G2X0RVRTWS1jjHM86GpoE84ha9gNrzVmgcyeoNcpYRcOnJ9xzXg22QBPirwuwJo3vAFI+IwaxLRz
vDbldeFcQJyQHRkrtLcuPlkE2Skf1BgGHoJGsI5gzNVcD1TK17DOLtvCM736R2k8SFL8siU9Pu8W
J23mNffum/sqS4n8w17lcvggwYtxOCJOOz7P4eAaKHMA83gaOCzJu4e1ae9uNLuR7dQvq15OmtzW
ctiEGdx6+FTFAcq0a7IVDq+IkPAdYWTw6QzbFgC0f38mcbhQYMbguISwtMm182BjNmG0GhotNiGF
Dx30n54QHoSdq5Yucg6cYrnGO1z714oGsu6cwI2hQEKe2C98E2p2Ds3T1nFKB83dr3dxB1i1vGSw
N69PUt6H+6t7RZwWOBaXL4XXxzlravUyAc5OZEXiqxk4QHL5i5sxSv2e4biWMr2BN4MRtl0Pck4V
n9CEljehp6a6KPOzHB+vmFTgDpwEx8OlZHiGcvSFh0+iKoegiofW15TLkQsclwo/hZkMAaxQI6Xz
SetYeunvbqsFpCE+11ksaY1yCKXu+RVyiQ/SjN1IYwIid5JcVwK1VoLBdszXliygdlXX1kANP5Jt
i1kHOOiXVTaDpmZGuA4etndi9HkxtkVGgv1AGSC0bwxbH1G73NakB6CLjpT1sMGvdcG1YhfoG4Ch
CdAJjLAGCpA+Ye1JzuNYYfQY9nFnHuceFxCkkBXUNxr76dAgDV/AfVKjfmOnFTs9zUNXD8i7ihOq
jDJSHCIgNQE3qqTc8iFRsOf262dnWTJb7jmWQ+Gmo5rixMEupLBvXcTwbybHw0v7PWBZYV02JFR/
6//ImFzUCxz67YgfYxYfiIhdJKMTLl0cfIoLdGutITxhBnEIIUeTuJ2/uDNZDl85XM3dfpBm2gfV
43gedBGyubXp4l7ZYg97elxJB1zlszXsLLcrhMeNNDT74BeLuNl4Qg6vF1suNBEX1wlBJdrVZHRk
ZtOKckz0MtnftQKjn4G665c6tYxTW6MOXk20cInOFDI19hT9QyqPWkQnr6iFR0/MFUaOFpAxPMxM
/SAyL9Q4/dV73ULPNZAZxjrJNhja5crOQHpngRiS6WZ98yOs5u0dYlHaYZ5Bu/65moCwXTGgSXi1
1AZwHDqAFSUIFjBBISKFuSQfZP1s9Mq/hPgeje3UqHe+SdmwBNrBeiaYiFd6lJM3q5LbIVoNOYWZ
BdVwN0aoRutLfIGGIexJ3ReJKrckU2rRcZ9FKy9dAP+Ml1kuhi8MSMtqZoZRI+FbB/2vgFhCYSeL
QOlkb6/LtR9ZJr5YFzR/1nGJ3MJcAEKR83Ariq95s5oOW2j6++uEePGrs5w+JFNwTzgYvp2mp7G6
c2UxCIzW+z05iOOSo2CQCem7q/YM0qDmgHVorXE7uoM46B6pI9kAVzmmPdu+07PFbW6AssaZGY5G
lf/9S8441AX1zWMuV6BnVXw60ijDA0swI3e4rCaKKwJ883+PD23NoY8eDakb3SYBLeYCZfc+Bq2J
YdfESTaooPc0xY0fwn6q1mm7yppKycrxxpYBHCV/o/eKf7+FK+SprkLGo14gOrdGJLkWdjXJJMyH
JXVEMlzF5Raognbdg6Vuoz9OgygQ2X7i1ZcxqWN6jE8EhVGS5Hp7Vu+eU8B9HUkMVS0XmmvY/sld
XOHI5i3oZSFyH7z/jUqQp6i84W5oYF5AF9VfDL8TaaSgylzwjucH6dbX4DCSAW4oifKr15hkLn3r
/SKALj/LdrrrTXLpLwOwVLDFiUmYf0vz96UmGZuXwmkO/NrZB0aYsfQzYjIBvzlqxKUXHW5nhL6A
ZGxyRNIbwXsllVKBOEckL9B6m0dLAVkOUig12R88f5ahsaoX/wwREiyer3f/Rgq9Z8rQw2EiKOoa
7UZq6ctdYkXzQ1c/z0VlBUZvldMnQXjzwKqBYQqH0twdNRxjr4uZZP37L4apN1kXj//TCRxGlD38
nZrMLfkGSpL6Zr3Hk6IkYchnMovdn6VlqaU2F+MuEB+hjsvTMd2rKu/JYcXEPa2uK2pxo17FfBw1
5c1SH1pR8xVBjwmRfuZVsz62xjBEvVDe0E97Kp1UDQydRZkKjOGmK3TFc2dFEQFGVvKuWzp+OxyQ
uyfVwrBJe3+OXGhpzAZygOIizohj08HS9ySl+nNqhwYExJI9yeI4R6X0myV0VLn17g05arLmALDk
Of0Gzdg1hO80XcKg9FVhLpFYp3CD85Hce3uDTpOj9ugWTKb4fLPumOY25ZV63ufZRgI4cktgRAET
hohBZ2jazaqt9o1hXPG32a3K/FiMNMnCjM6Vdk9Xx9HUcavv29R5lMVMSo7qi7yIdY3gkKQLWEPF
3YEAfZWoIBUkvxlL8OoVyncIYedYTT4mhLv2TII3A2a/2kVb2wTEbPGpIzMwh4/WnFtmHAQEZaX5
rHNaCh5vn6pKYt9gs1LDSjOjv4oEbGktmtoBgsebdOrLiWBdY3QbqJcqCBzu4VjOPH4A28T9iSe7
lnk1V3XvpBTAEwzGDXPfjzDO96kIlrT/jggD5ae+jfjoUvznQqtxLHhCxVCKnUGK2Rgm0tXgftgF
XWHnIhunxEBjTlB8Hd8TtzSHtpTsT9eApnzDOlwmbca37NeZ6HxlDOLQyezCiWZA0cGuPd1BBeUN
9chEDoVvjLA+AnbYBilUF0PZTJEUCOchfhYfG5lzofi++JmoVrVigpIRQKuihN1nlUq9bLZFN8Am
m663KXq3haMVkxwOvH6MoYB8IhNnZ/H/g7eer+Jk6B3wk6wmTvU1bPsMIew1sLoY457oN4l47bw1
vfJihvOb1kH3wWqA6zWcZ2Ar/K9n4zZgJ+n9gjcrhDc4BxIKtTxjEYYb0lrCnJQaxfSY/VQIJ78z
OduDQysLesykLbY2zAWh3mnhVA5RKxASaP8+s7BcTQiDronNOtZGDqCXS0A+ih1FwOO8wCN0zqQg
wsZgdLzAKJp9Y5PulB3HAGyx1NIS9ttQ6k3iAgoyjHo8k1ah+j0rGG+OhLioLPE9aTM8A8crUJon
+GXdUyNKdmhw6ONCcpbYohx08hhjDS29cQTn8XSxTsrpTCNu56ifwNlsYPvOtJgRgW6413COrAB/
JRExn93vfzVbdvgINqtN9pkGwk57/aJIezOVw46VTLJJHsxjkh9i14RZ9/oYgycaILeHw1Bb2jAO
3QIvDeicwMqgnZRUsfeBYXHNlBi4U/P1/0UrkpXJPMSODmniWIcY2fTmS7RKdcmLDCaqo/Of9sPZ
gWPVxvSX2IiU7Dru/5mkEyiKqXseJilJxNtfzcVIVW/CTgZF/MnE6eFqQ0xzMnjVWIJlQaUyjmPz
nDeBtLjxQ04OruvFx/ddfILil+SlrEzU/RxGCXoULx6LeFBQTgEwSi3Zqf/ZSTbSvxr9ShdoCLzL
08ie3O9JG5yDoRAzrQlcv7blbMweXh8nNWuYX7d9bo3kjsojIa0XfmePj2I9TcgXju7ZyO/V8671
6tz71jekDELnXZDZWn2NxGoVLbF4QMxSG+cZytHEI8pPfO8EFstGT/IrTJXKDx3mmpFOeQE+QNhD
Tnr/Y6sL0a27CyUDYilWHhDySsQFQIN66neB/1WbAwADultzNLZFZ5Xwoaukq1mHMvSQV5KEtV+Z
uYMJPjambE45N2F4QB9S8T2uV6isOkYxzaf8nwB7Jijl/rO1l0Wus66aRs7v026oI2ZIJk0RGX4y
D0o8WP88NI3SyA+b187LHNcuAVG+AnDaMM2WIpgJTIfl337eRua+w/dJZSiWm9dXzDAsPBanGv11
tcWbMWHT4Aoa8iQV2OrLN/AuNFjBcahgZa8j6Evh7i81Q6vx0KEP2wWYSj9QR3gDbaXDaVZez7CD
kBud/GMvVGkE04yysHp9s5fK/+3/E1F0rZQbnwbucAP77Af0gQF3sXG+wY/PICkWb6rFXlNquYnD
B7AQWOMYWum8xALTPqpPvs3ECpi+W1jjmQfp6hfGNJcHDsa5Z+TZBJX0nVSp9GwZ3DHGPCr2Y+Je
gD2mH21C8XVoUwVgVX302Pd6rSHz6FwH6h9o1g1KYi3f+MZPHCrcwqgItN3OKFpUEjTO6wXLxZ/Z
fu+Cd7NLfvMi7L79aLnr1Ae1PWWvA8uBd/ujJYQJwL5y/2v4im3uS0OdltqlA797k2Cu1EYTQPBu
7ixOWm4FgEG5i7CF9yAf9XuX6ofItyIJkc92P8fJwtYsuCaS+Vg254UPwfsaPl0HdeVZfMbFGUqA
SiS8xZuLYXXPyZ0OWy2r1CJQiBUXItNryys11wglzTXY/WnybDUuHk95xVcxBnuHPGG7seC9yI9d
CGGzbwInmRATXXM/3rY3jbzHEt6uQLLhLfP5YyV7d1W4dUJs6a2vYdI3bNmp0A3O9gD5Z7aDgFVE
EBEHaTHsUZ4Aq5lZcda6D5050OehmpIEaw3UFBN93AMphwOxO8yUSrGe10q4ozn0RtYye8sl6GpO
6PAAgL6k9ZN7Ai8nNwmK5RVb2FAhQQtncfzUYkqVAde3PfsD+MFwvr22TBO7PwOGlNvvNkyqRP6L
Jm3ERrTmMDhnJDXUEcMPRzASepWBSxkxLWzVuNKP23xz/XtKFdfVuGzdh4FB+AD8a7wiIbL2Bdl1
0kdTzpjyQChmb1eQPM5V4olEoJjuUMhlHTFevXs4dXrHwD/KK6F3gZ6W2P26nBJqRg7jOxIsX651
bwL70JauJFksrRDwlx/pFJdxKsiGo6rBC5vVFS7CWAGpMsdAWOTOXpJFxfYymS8Mj7MR06/xMpTR
K850L4nAW+3WamvXNdtCSo/UcDAGRs5XzSKktAV4dCvNmoNzTLkla/FA+wUDI1QFezdCwEKeckWE
WF4D6Z75YfGUVaAOYK4KPTHQeVOd8SJcPG/yvk+n4a1thXYEQvkoohryzVRiO4kyyUJfwO4CY2aV
/lmCdpTDDJJlr7Yg3W9JVJ1FZmWHRbaqHmkoOOk6RbYbxGpuRJfgU9028tYtcWxqhSO1NH+ZVrgC
NzDm/BXG1kWHyDO2RYrwYD910S05InyxNd3F0yznLzLoFQFqOB3nVVmeRdaaOdSgubdX8BmArRos
u1pfcTRrG2jHgj5l376Dsg+klhI5GcwoBOPwQySqFTNXkcEOKEWu9aCTkQhJQ2oQR9LUgZgIEE9j
P+G4+wlxaiBGTC6A47K2GbyJh4yAKvloZARCNvNAVd7t2hISFXYmlAqt5wNr5UpDj+y4ud1n5Ais
x8tT0sBqG0+sFKoCpL/OEE/t00tmzh3JEajE7Pa02NQJSOd8EGZXyO7GadnsvPcRBDUGnRkIz5vM
neqSvMfASPZTw1UzZKMtTYeFcVydK17nU/ZTa95N+sCRHldPKKJ0nfeJii8yISMyMUeMyM0PnK1W
xKKdDwA6htuI1O1wjkvnUD1hc3G0+aw2tj1Yuh4QjZE7hzRk424+524fDyNtQwghRrBgARKSiiIB
Qcd4sKvn9o8XBz3GudhaT0EAoxdQ7qyq2iaU//kmZdFtmeafe8xsyBJhai0SlU2q3iBIvzh6L/nh
Cm/6jR4XUUuuj525tHrOqmY5jAMu3SXHnSXnE6EjHKCF2oNMfFbJGf5silJ1vvVYZP3Ic634I4iD
nqU62hZbl8WCDqYFNJZRl02AUbLwGJZXy9ZLX+zZj6e60uZIOaRXyZg8LDJTl0qcSAjEqb0KSI0I
iAqvD1wtP3hTt4FebLSd/J6ZRhAIAksMfy7aD0SMsUCnZ+gRv/4ToNzcRnY+t/z+KmPwQBraga/P
a7Lqb9CMCTfGKfJnzGrZ6aGrlOlVxj5RlY1iXjA5Ti/OpUup4eb9ILjVz3GN0H3o0BFx1C/nUT1Z
KZSJZ+8C4PElfPX44s2WSUSLZvHH4bLH5OVdTzCSDAigNpRb3VqDUpulSgu76hxT+wStqFCxoFDr
K8Ug5Sz/XKS9jZs5vuyEmECDjuK8a+ISiBqP80OtTtiarH65bj0TVQqJNdqArtHPr9aEOkEXp5T3
SSTwNkRHTGPFAz3kkSSYk9ePQq4CrwfkiTlBUOL7KldHWvRhuAXL6X9t9BBJD3aNn/jwk5osYIDx
vU/5P4G9jjTyk297G+qbMG5Phl7H4q8t/RNhovv/0ASoY9IgOBZKsTlYw/Y/4M25e5gUGPgbiNbc
Wv3slgnSrI9W37m7j92d6ymDAftbWOSLe30BVTmHxagpwwTDtScr8Ckylk5WaNqlsA6fvQHiqAnR
GTSsfb5L1InXQMIH+O/f6oC9hP2KVpQmHJ6HqnrCMo7/io0cSDyUYMPKt6fdJWbh4AiwcOlX2ybD
FSm6WsRFLcKv4Mx775QJba5cR9prG0qzBolr0g+W5abIz8tO0+oPJnBdMNBgFgTnn4ToL2fwJznw
AdKHjysyG0OLSklTo9t7VJzUd3OnGTjPK4/byGtXx7jg8DmAkB9NMi/y4DFWPtiCHe4m4hVEg028
SSii9GibZ5EsJLBqVMm6ELl01CdP4r2VA79YVj9o4FVnxcNyi5il+EeYClwKJvUprIdO9nrOH2V/
+u2plYoy4qT3XpzV/yw0pe6h8X7ECsX6PTj1yMJAn/q16OI1RuCnZviGajkvKmUyLI4dbmUNOh8W
4OHTE+K4E0YlmB/eT7zfMt6N504a3KzKlNIMtxWvGo8XVZqhXG+7kc8o8Yo4sCSo97ZRIt6ShcM4
CX2utZf1IxKDrM1y7SyuIWJgT/f3L8oMFk9lB7ft1AOK69cfM+VVWs21qImMFtdPoS1H2BxQ1o8/
JesxD5kpREvItgNc82EszddWYpUqmkMGZe+nb/ANBsX0m/x3XNAokPog9Sss77An6mt+Mldsu4XJ
gjCVT0U2jyIURxzvYJvR4fqJKedTfqu0QRKm3p4wQtRUoLTXZhTB1j0nU+Tnbqr2SLL6TYdzv0ij
wC+4b/iFiGuU4NOlOslwElCMwz5hD87R8Iq7+qOeTv4zPO3kB853Nd7ADUO1hFx7+SuAiLvfauJ6
KzAXBCVoKgj/bUkcmynMCX0Sy6XZkp3hMc1tIIMw18blnA0iPy+Bnnfluw3d0bJGeBbtbSvfmIb9
KjmpgKwtauU67DgCcjeOdHyx8QxE0UR/yC3am6wHbqRRUhsfwohMwNRlh8WBLq1R8Ulf4eFVmXFy
fE58RBbrL1UXUYAZiHyIMJK8qpRdekQ6ErdyeAFpeLfY/zUAiozsstN55z1FqSyPrCWs5xblI5MC
0/u2LsxBhiTvquES9yhMZW5GTJ6KencWCfw5+Dkacpem2adetjSioXs3bs5FJkIgo0HaJFE/oZAP
Lk0O53gfLx7hpc7ILxQtEr87ti7F59skC0Dkxf8SsVdh0F94lMXeKaSSyMd/qDjvS5KsGPDKxH37
CsV+qaI4IjTX54eiVzC6UO/8Apwx+qqifhxg+LCilK27K+dFOmUvkBuoT6ymMd1K54fy5RiKoMUS
VtJc9cHlnGXRDc2sQZNF/Z4UdZC8SKlpSMJkNSt803LlWOVQ85ihcxodxqL9NRSF17YQObHX20rK
4UH8oWpgS4n6df671BtfrqEXMJVY9vZhq3g8GNEMp0cI4A4qPKfTp4LVf6V04L0nwGV9mo7u4AUv
tsabyj6+jl1cK3R9Pq/C2ysu2hVb50emdWLbAI63xv50eVj2oX7bissCGp2AWuudnf4SQ9Dc4+yf
cXZXzvbhIXy9HWwm1xCApTMyzZhCOo8ddI7sY3N7OCyErsObuiVdyyHKR3raW0p7BIc1NWlygCag
CDIj1m6tbd57+uEVxn9JWZsrDtzexFeFObLJjF7hkQG/UiPlOf4Glp5g2bCHSyXqIViTKeHo44JO
j2pzmF+V78LJZBFCYOTjBtosky0+N4dilrLV/IS6YPo9dG4+c76sgCAT4mWHPuwmeCmRouDskjVr
2Sck0uBlQEfVMmf7WBL9SltRjaFKRrGwLjb5atTi5ckvmLEan2PyJSWeKKqxabC5jkPqHtPwwa3W
1dEqdpOkw2414Oxzxy2UTFOjXXEQtLKtlPu4Vxm/zqq9Rrx64FPwWtprLSyfnuXV655pOdRtiryn
PVNs+2k21QB6Y3ZQ3o6s7SrUewEjBKiG0CR+GeFape3NUdzXaTd+nfl5uFllyMJdeBFihHieOc7D
xwtoWourLjNsHk2qsGKOeQUihEOELlZANfLOtw/RSLzASTdaN1BxDdnn6U0cpDHxHx+akOLYvDtK
dNOhpV/UFCu358sVJBHm8jQvZpiyDc3lxk2x3h7UiIeKJz5fxL5jG5v1Mgmh5jjlQbn+ARdrJDkU
lmW3hoOB0hcMw/9JiyQSY+72iHrB3O621RZxtzugf5MquDTphGRF3nZqWDkNWZ9VbFcxJLRXIjmR
0PWj3ZIKbKg7KUnJ8E4dGfMjnZAqAVVpZ7xI16rjrmXL9jH1PqYInVXjzgX28wT6ijC0UYSq5bC2
10iv/aeXEcJ3JGC6eRVgvPGRmOd4ZP3CUNc3jZd8LZCLewnqIeKacQOxuvcCs0uaRuEP24GEzLHP
DkWMYZslrBILhQN003Z7Ztxp1NzuhPs16Uyn2ItonFf8rfKGu92qaIB5ReYjPFQhX3ErdZW+KlkM
wWuVE7+qDt15pupp/0XMMoXcWHQr8HEkuyn5dUadqtl6PxsiohbvB3UsG1W6iLVFFeg6gZzYzNPe
z4XHkk+O5YQDQCGrY5bbsW8rMUgTLs1L/HiDvjVbuq+4iRLIZpwmMBZIgY3dyt2KI01oHT4XgwyX
3T1foPg43RBp3WRQRZ5tnXFTvWOHHEZ7lgARn2Ez04dyKmjJ0sbc1+VrD9g8ceXWo+CUaQ6SXAkP
Mn2l0zYFZIo4Bc0imraYXHt19EbK9Arc4eK+6UJSGrUsBzObRybWHpcTDWs8bteQx0joetVbOKmd
4QaxBrbyx+J7OdkkXwFJeHtkLWvwagqqkTh0vpT0+uzRUM2ciplRGlKO3mRTfvJCPsVYU3RkA1pJ
QFsycRoA9AE+/CPECzboWtzDvi6pIX5WFlCHfRMCYkX/3ND6qb5AfK6mB02OLyV+E1qLzFQxHIt1
YzUJBjbFDkQ4mTr0jQnEd2ysgRrGa/ZLyTSLPwL8w2jmCkLH4jNfWrs21hWDZWflAFcn/9hAQ989
nYxo2hTI+DR6L2Sgg0GOaiqvdaF3x1FmPNNoObj2sODrBGDtTlYCXELdSrz0KhaZYW3vkaPjuNIs
c2fQR4TNaqvITvioYZVEs6IaVxijLtsKv5ylcoPfhwLwt/NpBUYRP/P8cKQTwDEE5Jp2+dPPzca4
+7medsS0f3yvB0uGuVFafgfrYunm/YqfigS19jfmvaoDpSw53VvqQUYZOHz+KPn/Cku3fGmMx3TV
Bj6QJWoGpF73PPeEhIKzdf4/BEb1XiHbgO0XAm3GY61k11B3OS4WIIXWmqjnrJaATDRvrtSvu78b
WaYz814ohVitq7cDWpk2PfJDZ1DKCsw0DXFNz+kgUno6CjU6b9hNrOdSV5YSNQUDJkqxvdr7HRHK
j/dRH5WBIaGV+Ak2DW/mibSv6xGkDL686iHbgP0WVWMudu+XDfbOpi4Bgm/2N9A1696xFyJVd46E
0CaZbV8yNdiw7aN9Gyp1BH8RThu8jWA3jWlb320Dts0vRCIEqCXZV377PCmtdun9LDwBSHAXrdRx
oYKrZVAJly+Y8OrXsC+fNdy+ZIiuWY7UqjRn43Gd8BtgGhnm8SF+Q89O5aWUhYrrUPez8dxPRV0B
grJhPe6kDTwerLbzDqnEp4xxVVSR+rvoHzGMtZR5r4zz3bybdUfwEjHtwOsXjIM1dRZ12TRLHGnt
qd+4xyxfC8LcSfTRHD8JjzOOT8S0OqGxKr+5h/BZUHOHkdFpBt/DIQiaSCgvjKd+L6h3L0toWBGc
tbwRHUQEu4aCSE2fpWkSzQWtSYch/9rvECofhTLJNU+0IDGG7KdDPQ4cSYNuKE9EgDkuwZYuHR9l
l7rHuejPTKCs2tKB+R4NNxhyxGFI4gJ3LLvv9s6oOHDT4JvTg4EMpYgR4gVQvGUFNT75xRADusG5
5ly8ksm11fGqe2Y03qMCalG9HW1vUwFVzIOzfrupE5bKeplRvjQ96O2SV+AaBg9+7tBUDA8bYh/B
D8WG0X00nvs8jnDOPzQHtNoPIkz41ILa0XeTKFWVTFM47UlYQsNPUOEmqgkby4sV85CgLNEiolwi
9eGw2FdytR0f7dbDsyg2w9pSyFyGnAom/0UcwmpHX0DXM8ptoGaR4B3iSYv9laicLjpLEiIxjpFc
qwOxDGeJPnC9Jsam2twQ9mY6uzjKG41NoQi4tga3/evpMmBASMcj8NjGA5MJHDhpphZPUOVz4Id4
9s3rqusFPlQc/xxbE5c7Re644hyAhCOzX5CkOSswwgVQ4lg2ga/04kIPOFTT2YQGG7RffK2ICfWF
kS8KLIi51vArlcnkJKSqNzs412q23usqXb5gmWMDES6ZMcf0O//0UO1v+MnezJt/ABNtQXJYn4ge
rWxUXd4vRZkhtQR8lSh8Gb6nI6J/7TUyZKMc/skEvX94AeIpvIFydf8PwGMKbT+gpOixVBZaWKuA
UwQsl1544X4M/I1HsJ+gc/FmBREpa2JioX9Sjw2gGHICGZobdwICYAza4chmP8hHN3cqsXJBeLpU
aizyl+x8KhPmwfU9AcEGM8rLV8kwvZbieWpPqJz+B/TcqMMMCfRM4oRcx/AfwwLzxB2Zo+ba9Pdp
mADtD8GkM+KsbgwidKDv4fuutUs/2Jo/+XC12V9XFdST4CEC6IOs3Xyojywvw2yiWjVcRghbum8/
NTGxFmlrjx30pwBoXg82HH8sLZHmW1Qx1SPCIRWvmfBkvNTRbncd82jS3ooPXhPUiCBM7VfIZE/2
lHcWnyyEht9zniGROkYLcket0dAkSkg2j6ZbM41TogqDsdG0n+y3EaXD/kvjqgSk7ebIlOBJfXrE
XrIQJMLEDLWIapRpImNg8bpdKNVkgR7OIJrdq0/dFuqRtStJKj9PL9661EYTlFdhBFcM7LsxI4wX
nhtkHVw7L8w6xQfcu+FFDjDrBNJIqGJOcta2W2mA/ZxFEW+Luru2plueTSVzhhNolLbzvPskfAIg
hubSAxkwRfcULsTAo4dU5KBX0lD8kNmc0n5oSvk5uYpK23kJEUOwBvQ1ojr36zsW1C5/6LxNO23m
au5ey5G1+mEMh3CV3IbcEH706+NVdfP3wxnP7SQRfLwEgVsAgIb446CPFdcZLiZtAv5M+5Is0Joe
HLLHrhqy2d5+u9Iz2pzveCriXOjlcevIGcb4oUn1A0a89vv5RpCGHU2NR+QdSiibweLcXQXqnoY+
kyZxTupKUTYqFvFjmLHS9uppzJytWuzTY5yaRNsAb+KX4MJLobazmv8l0JcKe6/EgmNYulOj0SHW
aqp617uQWRbMk9LPpKgj4LHWRNbmmX+rLfyz+LcCAzvJ3VjcQh2VxhopKND5JKXpgnSOzijC77yD
i1Xzp87vqZ+0MkTu420WMZzf7pMPApDRZYIvFsZbCjQz7eqpAjmKq9uUav4WM//h/LXNwF3NtOVO
rBYok3IAqP+P4yqwS13uL9KSXBqNrRK4aoxjiUPvAEARX3EAJ/uy9fqjvbaT6YjkYg05OICLBjDh
7wYS42YaZemA3/wM6BZy+V0FLvr4ZC+urdr8ysZCoVmhFlAWwhlTWbuloVKoAkVEPgNGE2oTd/zb
WMQ2BqPilkV6IpTDg58Wr/hYQyn0dfrRFwH4bQlUlnQeO/Lxt6etmPaA/d8GiFFzcOjaYIR64CJC
mhAjWx1w7Dq1qs3MMtwwtoxgYq9m9mOMNgQr9P3S+VHGJ/BXp3SASEPLCayAgjg1Ls3rITRvPRx0
Z/zZXhAzvo8gfguJzcoGoYy4NwcWCyzfZ6pvQSB0Pyq0cmbWwVXRpUckNVOsngfAVBRNw+PdfyoH
KXn/c0IOGfjiBIosK2ATky9KcVnsuTDda2lHu4TNqMBynWEoCcDze90+3PGtkcIylv//DeYrHEZP
nLhBUHwv7gqeTLwnge6gjgdWhtZyGIoar2VkdwR2tQoKIdYwoQzFHj8xMidLhbuQXQ9bS6Ey1b+3
TO7caOJrkGpVXkQQa4zfaJseNxdKTNR7mbu/e+q0oGEmZMDbJ53gMIzDNFld7SZeFnBG9TUlLiAb
ASSpFwmVBlptrfbFt7+bFmwZ7vtAWbMIm6X44ZnAzihTpueXQOmyeKhZp9GPqaHG1JcGM43PWBo3
VcJZm0I944PcRL5WmCf9E6NegunWx2kq1fg9NEeKKtmlr1sx05HQjwmF1z/XJz2Dxqj5FS4ONj7S
y1a3BJvHKNDo88siNLeVDD8KEL+2w6gyYzJgf8shLbXfjiDydK1vk9YpMC5zIM5yWDQ97bitaWdf
9idmjyA0+j4hXb3WtkZIUiR8BFqNStydo2+1OckIemgbiFTWBMDD215iyna4/4niLepIPMESgiZA
i0NOI2W4xdW/xJ7ppqkH4/FbJyP9Y1mF6wRVls0O3EJ51Qzi9Wr9ITU5DB2p4HQ7RV8/Ejk1TGE9
PILRq9Tt6JtTd3X1vHNtT6LJo0CXMp1jwPhnMxU3k1ck6stgnMLLD1YuL85nOP/03OtT+EI85a1t
raUlpltQo8Q1S9s3Z+25AxSArOg2OZ/uNs/+mFrYFOTq1VkDeLt0EXXLG40UUshRliSpnT2mzQHR
oRhJaS6nUyJxbEK4A/klVm9oJt5SiGL/H27K8GzUXTAGs1Qw6NryhBRUEXpiUvx0uVM+7nmUbB+q
tKZEPl6iJi548mrx5dYWDuBcCFfwNuDDd87PLu1ceKSdSc9hXTpNexP2MvlYksBswy3yUq6cDm3y
DBSWqi+9uH3irT3zV8c/AeLICD88OjhZXCit5Kg1QRS9dZAE5DvR1XYnfsP0dDxasR8+hHb4Bgkw
4X24IawT7p9o5Mf/4/vszcajp6AVX/+2tcrVMNojxcA/Vtv7XfVHLp9Ct3NAMRxjC/5NvDGup2ZP
0KRctzf6m4F1ewOp7tRierTnBBdv2/C0ofDIhjqFRLVWj2qlqPV6nb6TyVroASE9zH7jVDR/4jqV
u7yJMd/K/lfTG7Oln3QhQSZRAgRycc5sG+USVdn6i1TumjEe7nk5G7mSBIXhq3ZR7zXBUeWxbcGo
chV1EFisxL8YY4Kmdq+eO2HPRiIufvqlo6q8va0wolBNTeGTc4HNfSuSr4lFwJ5OBY2eAlth/CZm
GFOXEeH0BtVa1e1rOceNMZCMD+bT/HMzROo/cDfYkstgRPM7oDha44ydHvxLTSuJKM0xljIswmr9
rIs0bc/BpMUD8xJ8uezAErsC9Zgtdv0zmpIRdVDU8QPkzTYLjtyjT7noJRo0MjuehzfxdO75Lng9
dtoxOnKsySGj5AXkBjy2BxHvmMr7pLcE7aHEXGGxhjMe/DUqhEiUwVxSCvC+mybrtdbXglMRqgZf
0IEUO2MbxV2dWkiYuimA036c6J49T6mLpIqYxmbNjFguwUt/7yuEPuJomkFEgkrWBNoZIIpU0vuR
1t/kW3NhJk38jl3czpR3kyBQPTEfW/kApqxftKm4d94YjU1ZCHRBCSrxPccEnBeX7G0VyZj8cFpV
Vr4KB0Q68hgNVv59bR9TJbuiMZK9gKoPlAHtOoV/fTfEggsvoS60OZxDlZPt531rSY54ZvCgp3gZ
0XShclOvP2W11MOPeaInUHnseoBFv+3jphyFaTr3xlmUa/Onc0o7n3a+f67S6T7u/JIiEgf4FSzl
1gZD/g8dsZgGpvxitPcTDecuYuP+ehF1KeU7MqC+hpSdeBnGF0c2Gq+OxJZMqkOh/72j1Ad/M+64
vdblzrD9/BML/NRqP3hItXDC73aDMCfbVmC8wjWtFR35QTF53euYPrEcqh/HnE/jWRAThrtFSZE3
8opYpyb0FtUSdh/BqvVqsdtrOEJSdxEtQQDCrik4kXPBMzZqjJzZKr/Txzs7EyctSowkjL6MBPNm
+nUGMWiclhf8Zs6UGsAb478oWj53qk+Q5NkYMUQnfwE+PK3aiNVPMey1X2nJIJ8G66Krj+zjaWXb
jeNIgbwJp+VYgjjTZlyLaYCVNNkv62Y73+x7TXk4eXLW5P+FIM2LsWmlVJJukRHlT9IKKaymAFSe
RnekS6/mp6G2bBdI2sdBpOmwCdfFOoffAnGbcxwxQK+4ROArtZPWJ2FBUvvAXCHy0SS0PkoxMpFA
NqqiiZ2/AI+Z4/inYbVGS+uy5MF/CKkHD2zGyUOGv5BGPO4bvuE0iz6bVnpfzgF57s27E6yeUZW1
nb6BuXccDIai4mDjVdQKPCFS8b/4SsxKk66UF1zzgluT/nIRNV77W8SppnGvpVVflde7t43pnN91
cQCsuQ3B30/xpSw0pMsTRq3VqkaK8xbwG28N7XHhBlWizg3/MSfY3a6Y2dtOESpFgFuUCO/Dx5iS
xC4MCoZ1QCt/yZ31YON1ym7xbTiPO/AVmYmrHvO9fOcO7IQHr/23EB/pf1buNHZkyfL2LwQIBCzL
NeGe3E5lr0SDHo3z/qTNAys8sDBGVM2zrJGOcKrCUtqWCEkpeXvgQChgx79Lp8wyg+OyBsoVEJhH
fB+buPejwFw3y7GpyviVvvtqEXgg95vbjXRyNQEPxUoV9/nlcMdhZT1OypGoWV9onbc99RLcEBb/
pJPulc5QhPQwDaenhjlVDfiFzSmFop6oxlquW7kDV1aeypwU3BZ1nxLh280Zv6dfCjfIUotN1iUo
X+0Ywt40WXHqDrrfpi/yzy2zGCKJ2K4j3ez0NWKfHSYT3IHmYIhTMnQGyYRNNd+bVMRMhinqQWxc
MwzRSEYDzMknLDZA5e0bZ8Uo9pz/pVJFKAlfp/ZvJQz8F42N8Hy2JnkaY//tyd7QkoreIUwOk8My
QXDUFizjHoApCDoLTvanC7/YpUOs3D896Foh8ZlMuTl4tVKQsttsQDKjNrQPxZXQ9howMr8jEZoP
QLrrb8uinzTFXNkKc3fpnjee47FIKdBPJ8IQ0SnEV1CsRbf+EiKIeteOedKaW5dT/tqHVq4zLJIL
9y++qU+Giuz8uWR+q4e/I7nvhR2XXi5fjrh+pj4+HHwDa9z4KZV5tCbrOcomQzUFcKKOe+iTbILc
Snrt9MLqr/ys7n43jtOgF1XcppiqbdvNxF/en02s6oS4b2IBtNBr0J7R4IQAFxn4Yay4kGIC9dOC
QdBXobPPEjeQyT65KuWBLW7/etvxVyT/37GXqQo9ycEM/kTWnetz2XUF22dKDCP85GaY0O33gWx9
C1NKdKSTeoN4DkQtNbmk3C2CT8G/G1AtDVDpvE/20JW22pZcFGy/W/JUrXc/btA8tSftbR0Da0aM
9X5qzvELo+/zbIJ2wsNtNkKiYX5EWxUCCSWFbkkz+CHjSVjL3FSlbci0t0aoEhPlklp4uNt9IAnS
QWCUBgTg04WiWGfZ5fn5G2/+Z278kuMm53A4hgsYrVZrsgW4u2DMnM5tMbwUye2Wz8slF7tme1YO
cEMRDyAQsiAs5nRh9+f71puQYPDGgXojZJQ/BpLkqDNZAS1AMAdgPANjq5stbBCVEUFQlaIBb0a/
0P9SX0Rm3v2dQjnxoOU6iA3vH9zcXUk/bs6nq7Hi1Poci4jJuFgsACd7ihAk9D7xShQ6+Ig+1YyL
EdYiGbaNezH6nu5l7AQcKtPPR24Nz7pmOMo1twALOa5bkxgFr70QAQBpHV8Um4X4wafv/V9ioRDq
Ln8PNJdDPQtt2HkJTL9UGcgM7Ks09toA2DKWu6kVeGG8m47wUvXm03HW+1TxjKEakNoSWD4BUDRY
5n2asNRqNtNhQEhRNGwFyxOsvjlE+PrdzYlwXnhxMEUuGdpqOrkJlp3zEeRbmiQVWbsxBrixf0/f
0ZlFXE0j0hK/hNSZaTxlmIvs84vjQIOreIZJUlTsFTkdQWDSz0hOnX1ALvl8EbU9np8pn7KLjz+E
n/acZCmQvrJftM8VKt4pX2IqDUpHbSDVCPl/mtOaR5+NTApHbJOvnu9ZJLqxFxl0ZwI+1KZ2VLZW
khHnMgSzJVJI4JhOiGwl0H6tMjNTW/WCRAOoxuDb3nw6K2/zuzQdbQqPbUI3I/w8/tY1LcGHXjUw
pmd8H/8k3uURDfG6+98nLOkpFvuzvQZKV+IGYJlwcY82FcrwIIasnaxINjfgmw7Ddd0Pil0B6apG
6U1ax57GNoDi65qxgVH86UTu1wWqQ34/ssyOIsKp6dW0BCJjB+sZql1VeG8Cwl2tK98UaySDGGVe
PhTG4XlWEDQ8zFGaW3FInHjr6eS5YmYjnBnhiMsRYBIL8NsyuVg/LhH3STbKvAUYj9nWGtAVBJEe
oAPaCRefxZ3rj4Ou0UEPBKs9g0gvl8S53/N6fAzk4sGP+fq6VWFINtv2tbPWSh9ZjiGoHjYlwmSi
+h1EUCHI/elNQjb6txxClwAESYF+vWZDCXjg7G8v670e76/FqDLjsP3FpV6Ljy2AsmtIP/8ZpUy4
NvHpVHYlUqPFsJ+rza+BPYvdfE3fWxfQcv3+qRu0K3DfncoXZGFdfYMlmiq/lOH93mwDLp9k5+gE
wH889rIUfsOYLGkhSBB/RI82tPnNjscg9Hd4kZo6t6oUvIE3DOHO37unq2gT+Vn0MDqT0orDmM6N
nWE2f/diifhEKpYaW/jXeckG6VmVs2gUlJggvHUpoR6+ZZ1+HNBwgpF9NX1M7DA085800lTl2pKl
nUt5rPAc4DCwc8uBLOFfIieSSRsssxyf7UCoF/+220YL/W1yljgSkJMZRtM/Si/Ta89MLdrlrpRN
KVr69FR7OphvHOZ4lHlY840YSdApiiOvbif7lPMa45QJDVar0lyL70bisCu0Jab71TrMzWc6YEl3
I+LQv2YlP1l2h8mgHlsq8BMptEvdBnGCH/11NHdn+wwkgEXQxoygeKbvFWu+JXfUyXewtuYCyBpf
iPewjsKCLEjX9B6HvoLv1WyeicbshXrCN0BiaStapkRM5LY6TrKCu0dXIyO+UzWiCIEIVMrn0Azf
57+OWCi6cPfH8G4hbpO0xPWaADlPORmiJNbn85/O8lvU+tgKLNOOkvIZWRX9vcFjrHkbOkx8eWOy
KzbIbSI67UCFnpvr7ArIYnqM9UeVpTYybBjRzyguOZAFx9mloXR9GpbYNF6CYZWenimSBAvXwt3e
DZj1Vr4QPrg/hcC9XHuvVY06RNKXJzkHLjpWe4Ij+vqdDYLmYhtTocDFr6vhIrweNzG7xUxgpi0X
muSxCuSHpuI/ky6n8bMBV7AWdmjSWgWUs2ZMexH6nbITzepIjUh165BSLGrMAY5L6WbKK41h+TUN
Nd/g8e/cnH/ANkxnbl+eM+bjPg0QSwJKk3edY80jxKzLNzPgqe+ajbpPHXdlZieoQCH1fJ/9dXbR
ZxH/52FFT+iqljfQNtUcRM4q2eMr3NRNNF4Y0l4iF85Cd32QGRXhKftGg+2NI8nfXxYRhZC1R+99
J6/A6zFepp2DNWbZwjeGKtRQxZUETvNHZr4nYOpeCBqt6inoKRYadVrGf+MBs7Zas7iTtJKBBlwi
R5sg971YCgaMV1KsfWvH+6GuygYurpHsQOjeLd0qlceejY0SV4/HBbyEPDYLVZ+S+oOJeSBwsjmb
OAUERqoHnfg/6LneKhWfl7/Z9CvVL6Pmj3e355bGlFwOeiIdlPdrq2pTPLPI5mbP/qQ5+zGSUFrR
g9HgllwmVNh1Efl7MhEZ9bqBEn4R4t6ufHVXj5nstoFnSfm8GHBDP+KDCJ3dw04W83jjAq6Hazys
rmQRXf2WGMutgGpQ0u5OZH93Ph4siin2lhTpKfKXlQ+dCNcNr3VJPF5QcocGRy/kA3yNXpiJxV3n
AtpNX708ZHCSm1D4tWFa8xIb2tib+qqUPCbz/kn8WLIq4Ub0d1AHfXeUGoyqoYrVrRdjwB4RuQWA
epF9hw9x/f2N9Eih2gvrjr4vvTmQOdpjaOWH+w+PsaT1DPLDL+0oGqymNB+dxqouj78oWV1r3/bY
P7guo1eviz0pdtwFA+J7dO55dG5JdrXL21gn9OnakyPWxcAiUFtNjud5/ebWSQC2pI6UeUxBOCDf
AeIFeVkwJBAzKAqdmJxU0SHzMY6B668g0/XUspQpAN2DHUduIhDroi1GuX5eUtNf/UaFH3BPeV5h
GSPkn9obHPAgGoyqZPAiPpfW7Wv8wAllsNF8paDeQdfCYyrp2B/jnHjSv5jRNsyVAYxYNWoKdw9i
K8qjUqCVw2qUMpOfUv99VyqAQKtzdN3OSm3fd4lRbuuAOkGGaXJXVActdJEb4jcrkzFgA7zzJkGv
mAFTDNa+rSGZ+GVngEqcuZbS947XvL2zci8V76sw0cqn82dCRetbxmKIby4LZU8QFUfXqSVlE181
p4887xzySMxrM63i0rVojyN4qjEbDcaDapRTlqTa4Dhc6YSH9E3UR7pfd5b5+Kyh/h1k5SDzck3x
mJVxQlE3lsHJVTQ3O9xHSdzdH6nST1Lp36ZL8WR+lG/SxbdIBFN0hiKYlLoPHh3GchpQKh29HP9E
zAD5iY1oy4EKz/5ZjYoQrn6m0mGaN+MNX9cJIwGFlECdWamxRggNagJ3+FYZClLg7BEZlg9NiAyj
DPwTFtd8Dgx2PmrfvUkd2pEMWqfz9Jjn98GVzKS5whQjNmbDa3gwaPMTRCncZ/QicaKc8C4LDyi4
gJWdUDSxD01a7NgyDy+Qh6A9VaV36vMHFx6GDZDoAonddsioi+uIfeDnM6TzRsB9wBmIkqchOLtk
2kin18A26l4RhRzqNQ+xYzfRO7TAOeMmHcymGyAHrAUY2zpMm11CDBoxCBa5VoQf3m6BmXzpT+zI
C8scpDoDs1xdMneTce+mkYVtAVWRBEuS4tDNLeMIaeW8UEnhlyUNVggkj1wpVDwzaxHKvEUbUgzb
PRTkdwqNRRbnDUdy5W+wzDPEqbL/KMfuXz9+PEKxsuL40Z9f9FYj8V9UpRs0cbWTvqrkMp7Z1pbj
5gJm92FyHUi0iS4LIiie4HQjubEzPTXkeXfvUPszF+IU3K0kGL0kHpHg/HeEXlG7esHW2ciWfqQY
sqbUxx3H7RviCPKmTxhDGQnbUOeUSNY7SfE06vgA9FAEUPNL8PuolNvEs3L24PMBg/kruFBY4kId
YiT1klHjvm+IDR46cqSKK/QyOi1JfBPn2CI75reUcoPEN5tAqonMKgPggS84XEe2sg5tSq7hEqFJ
+IgRKqNM+EJnxiDb1P40zI/9DICPnTDt7QdChzP6ikwONJJhQPWcKIrSo8Ie93Uot5cgHRg21Bc2
nOHaqHVR2p3On+h9n3HMojxarqqsqK60h9nKJTXq4cQumHCEYSGIEobCyFJCwn1PW1FUAyzyTKru
vCQw5ZF7YkYahRhQ0wkzID3s+Yrsz+C4Qm/cdSucsKgFogeeoEGDfOQLHUkS9IZG/LaT4rReulQS
e5zaQ6FQBVl3Gz25jpvUAE8plAJawEOhBn6Krgyo9pSLY7K6bGdh10eyilwvYplNHQ9VSibOA8Vk
+PW/Cg8fQ5ossgy2m1HlJm1373BZ2tpHF6PeVYP4cWv5+OiHGsqXoVPBKpPjUTSJT/QeJX+2TXgj
1em28ncwvnPOEp18DSa50lXuQ21dYgmB6ikdv1rsv4VeUn4VwB057ZVqV36/aueeweWK6SKTKhLw
Cvp14UW5+CU76RqTtafndlaT5PfyYS6bKB6dPjo6CVv17I0rAMmSx5MekBNUyvU7Q9QUaYdwHqDd
DmISaa/sqlSaZLOZowueUSDlJd130V0IZHJIUkflA0ddFQrXCRiX54aXXdaHnC11atavrhkS54cZ
OdZr4gw/GlhkTbj5AbgDKqVBcbD7mc//20zho/vRZrtHqDbekygc0+/L1WVAbLGcC13E8S7fs0+d
EUTokpJm8lRC/ijVy6X+4YLCWobk6XC3VsQT6p70tovlHXNTtaC+sbibLlxJxbgKPQWnWS+eX/y1
Oe8LbhwbE5hs5P+cft2bc0YkcaEqH/vxTkVA2VIgXeBaFC5abFERckwZk6XljG4x8lvDlDKHhFol
CJ8x99rO7UJwnzMpLvSKq2UwGxCxtqRCXmYAu4gH2Q7LPT90cRkRa8M73CttQtbcDiQGT+ZjEBfA
uSa7k8Int7djIbcwljDJQP/rkD/hSMJ4Qm1qxQ1ar0AkZnejm8DtCUkm4aoN5qHRYdab3yjNPd0G
1xDGBPngAoGpDgUDbBpRIII/9bYGwSzZdCFR/bbKvXujEoFrXby98Ok19HczS8WYOKDZi+/5nIFL
jUq07KeCl9Xeh73oIYPgVOwJxhnE4Kr3aD02TrEEk5/VkG6Q6JTueujcDpQRs0ZN2FDQoGsDUGbm
RzwB4fpn65CYujio6r0mT+D5UiqAMNq2OVYOjwfJ7+hEAeS96TJ1KBVWMiXBDM7OclA2XIOjZk8H
woHZoclDZCT31hP2URq4nRz66ynq6cHTjFAe7zr+cbuKu0eu/IQzATtkDBIYlq75PrQFIC2QgUOH
pVenWVK3ldj9nhUcf+KnD0Spgim2e4LQI3Y9ohUAHPmVWoc4itAWrqbLfZRzbWAQ7+BsHxKgC6hP
NPLh3jUaPJfLpP0fJ2kjVzuKCraO2y28vkdIdHPzfwIqdDYXmgAy3AU0FEhmWq/bWtOhtRqPJrWw
zVEfdTufVK5hguJI04eQghmvUpJwtc6vp64ouxH/0PAhwPNCAsaBwmMCII+idohfNA4b9HgT5rTz
CaaSt9OxtMUzXOcywVWnaPkdoX2aDKO/6/JcPtEhLTk3ZYGp6SpiopB/ORrBPSdrmWqY5aa/BJTO
RoBys4pa0NPKCxmuPu8DlvKAdLQe5etpE/TRYaAlWNtksVON+b9pRD71VJvZVFug8lkdaYR6h5Nj
jVSk4RY6bU3D0AxDp1tGvHb8DNi/TEiy51pURx8qP9mxNIiB0IP8yDwFWrAxxRunrlnY+h+/7NC6
p96QuLSpNZYas5Nafoq1iVShToycN3Mz4uCKF2ZWTn1/EwTlL1U+O713Bjjw64TUgU9VSoPbvZXl
vkrRo9a/MVEtTF3lGgp5cupvjCgqShqvYvZBtW5nRUbb4Fy7zHvTUgr/8nVKPoB6fCr6c9APqF56
dMyuL22+9mZMAmrY6UYrXzkfAWeuxPJtMroU/rJ6zxBOVz1I/c5j51JCc61cZG3mMegc5sBNIeuO
DsrxKRHW3RfDtNuAB5cQijUOnxgWBfSogRAcU2xVayGGuHWfw1d0HYQB7jwVj+XLLdU/HU75sigr
oikqnhP7lzY7ghqyCNtB3JkDRcWXLEq++prKewFRLNE7f0xzabGP1R9ayUFgVDYoINvvguF84psj
014U/POu1+QA0K4nLhwkDBzRRSVlukKoCGicjsSqDpNZlkW8sIIMmUlQRlO2CEAjqO9u6UVIFBO6
8SdiUEmFU2zjjPqMbKepWFZA1O+p2J/g+Y0gGbpB6fobS+eLNjCaZSa458a2K+7H+gwthH4YJBjI
KTXIC3CuCT9hLUK/9f0+Lyb2Yr7mStD8WnfUb0cYMykbI9oq3rNl2wV9kiwzB/MFffwnz+VrF8zd
7NCKAWjURxQ5+GdmpYwYipi3wi03VyZVqHh3fqo8eYsJQzQ/8QrbFGVtriuG4aWDF9YRQEs3I47G
vcnvLPdOCK1+iBJgcNKlwUxdmSExSjK7rOsK2375nNMHXBXhuN0MU9Ja17SazSBHt8CwUtqW/vAy
tMFHwYp3lYlxzIPpN81PAJ8eTlkPir8p8ohO5mWAxPh38yYzzzoH84KjbXqfFq30DxJx6EB1rUPy
AS06/NCtIbSHtlTfS5Vs0j6se6hnotOOE+y1bjTsjfvbMl/mR9dbyZ5FCHi703e5yRjgcJig8O2B
ONJQ+7WgAqZRGlRzfDX+f7ZBu6VMMEDmHCB/Z0utKsa5bj4uZND6pjOpSJ8biphua3mMxjprBREw
BaqhPBsmX4uvYROdiRWJm0ndVqHFYDlPzp9SBqmZDPEsLGFEIH26Q9sO5VD2R6YL52ZF1pIVO2jU
tbx6ckhO4GEYtTh/oxebk/lZRTUjz1VTRytqM7qJIVtt2nWweUNcrqPIuIxxcXTIdmkChjRtHo6a
5hzs7jt8Mz+n3tzPHW5mvXH5A/8B2+sezg5qsW8+2lces1cJ7M2T6Cpz/noOu9/HN+D9qvdEI+nc
IEtze0YuMmoto9brV0Qu4F1Cdu95Wc3Hsa6DFDc2UqEpuLDN1MgunjK0d09tT9/GA0GuBQIkdbW3
fWILFxu4OqyPF5kK8ZfS+iyw59j2S4tA7aXtCBTgmwyQcRO/HIeyOXl05BwK3Bk9LIFZ+KzP0TaH
ivoRDrJ0gdZJPSXUfxrgn4W466pQN1BE2rbqJzz38jGH8mJ698jqd0ZZ5JkUYLRA4BDlVYRF2Ki9
qS5OS6+RkkdgDf7OZ0tY5htsDX+2pLyn2njX97df4pcuuX1y5x/XH1KQF17yIVtwAV3FnQz46uOj
7e551LJZQPE6J9eFQE/YLqwVCCysB26hdGzfAAgLTqlSkUMCEemitWXEbkrFOeh63L6ihbedBbmm
+Ct2WWCWQI9pC0CDqHQcyLcbmmyOEDKkSx4moZZZl/loEH86RUH3rSJqZEQJvlUVUc/j1xfEitxO
3GbISdmyxy2DLeJsIShLVLtqiIHCVVmLr60xwmSvLEZ/OO/oVooTcdoFSGR6LlcwmO/86hjWWERu
tnXyzlvvWmyCwJGYRx4rlKBh0doUTlcJP1TbPCNmbXUFii0jtSREfw8Tp3bLIUt7ASCc32WN2B15
fuO8spXkslalT0a5AEHMPMKSiicK8rH0v/YKYNlfvd+gKFq2UJT95+XZyqTPo57bIaPpm5pUDrAd
Hc1R+KA0PQUs5Lfi4NJtNNw+QTmL+R6esXFJicJVZNqhZuUXO8ZMdrSxv2NBakw7emEYTfM4UkMV
HxbX/aRvGsLcWTyysoEDHphv7AycBP9aBbJvesTMkypbV2p0Z0mvgmPMUB8n0+CwajaZtTDDqPlY
+FKGLey5V9yzrxi7NXNMZQsmaoVDmxxBEhZsCji5zYzcclR+AUq3WU9eJN04y6/oVHdx+eD4pOos
Lwlbj/1F/WjK6+dR4+PGApJdO90lz7FYbUTmbyXjoendB8ErbwxpGe84JPi31aFn54plcWrLGv9t
GRKQvdpu2KdyVvIvhoWb5vH8WHwElzpN156D6mnaARgXcpaxdnJHJc1uwLbRamg/yJ8xZr5h+B2X
Weov3yYWDkw7uMmudVGoR5z4ZCvCnQ1I1jvR43jKKbcq0Q8ZS4w6RyQOXqRKGrcejGXlXtDBo0nE
NfRZkULmb5w2eUA8PWp4mBg7nE1Kb5aDyl5cOkwSnBaCI+SA5+h1x+JWHcikFteyb+jbSWKiB2wY
8KlxFbqKOU9LeXK+WZxYbF9IkgV9Rj73bVrX7G6L9P3zY3PDgAB9O+lh7Wop7aLi8FasAX+Vsmkw
6S3utuKcoF9ed8HlDGpzKDd9V2SvFnet2KDA0w6MSo5naUC/MQ2kApHJxlpAVAPhZB4S6ihEC37e
5ihFwgf+O2QcuHaA9TXuRMqADGmMsikDoi0pDPB/hZrFIyfNIVByGxx8OZYE/6akvH/d6Yim8AWG
Hr+fFu9b/dimZem+rPNLtkb1UahisLG6wNY5sMjBFFAK4sY84VIQpXfilWOPm7vfyK1bz51m+BKa
d/Y4JRckqNu/y/9KSOPca0N9q8ZxcRywCxM/01HXst2ewtifIwafXv85V8b2a7VXASSNZrN19rit
PS7o2+2HKhhA7tnE+Y+Qen8WPnTw8ZJHTSARwM+mz7mpS6zLg0wU5EpkhShKbq87HIRXciteIxs2
ennpLuFSk8PtubQVl5s/0XXakNb4jsO/ggQIXktt9SXbzOaHlr9fSclgC8UiKZKMTdkC/wfTBvzy
L95/hrhRLCxYbSPv5mAUjepxP0EvOR/a97m52TAp5AmucAKo1UtZb8a2n9i0eU3VksydpXUVC6tq
+o34zIHO6icbA8iG/fzqC4v8dkKsiYs1Jevxf7szANABrTsoHl2/NPuS/BU/Ln7uaMW2IRMKvWI1
UENA+TYTZ+ZQksvAn/jpN6csQzYavyp7lwogzr/tZDq5ngDsSOMPhFdSLrOuMvb+k0wsfsJmCzjZ
fd1vbl4qXJhkTsq6CBnBb+Q2qryTamSXKcygZsuDvRxwqO5ZMAXZbQJ1eR85omn2+8EhmyP5TI3Z
CIV55LkGwhk5D6bfzIhx8Wpb1GDP2RfFPuORbAs4EcGCr1WUlGV+5zu3GfTTuZqkGoyuaFZDWarv
6aqSinSV/RCK72s3RntgoaCnB/bASJYM+MUf1QTHlSlUuNmRudDDgcUuVR6gqa8uddCqiijhoCNx
uQoGSwE3lX5V/nfkGmumMQ5FF8T5XoQWriv9r2Mym6TjZnl2IgRlgd1UGzFpAehwmpmbUVR8pmYc
Kny1mFjjhRr7igFwla1k8oGaM1liJM98cNvC+QdLoXzoN7iSPk4Et6l1ADdSlzvY0AYXdY56kAcx
RPeZfoWHiP4Q9YMsSG3JkBzKRz5vql7JC7N5PCV5H+srQuut0AaNraCaaFOLaUJCdCoPj7tcd++t
ARbt49Fs2OFpq2IZHWwsIYJ6Kjro/Yhvqdr7eZvkK1+Zc/B+kiDcCGaXea9Ch6N8YazLUupM4txp
ISxZTcR1Tuvgki3CqN6m0pE4HAn4yglj5q8LWrcSMtHAhwLifonHzJ4ZTIJaG/399syk+vu0LnFf
nNgSsB40nV82V6vMAtzUuYTmokHykw8jJlTZZ6HcmzAgDsG+Sl0bXeLvnSRjl4c8EuVuYhIyqVZi
OYyLEVYfciaSBT53WYo25FkwPXo4vgbGeA88QEdVnGnK3F8tybIogNe8NCNzbcAmGy+k0Xvr0lN0
9O0vDb/LYMHOoaY7N6yV6R55bZ3LelwOjWj1DxBnQrIoC2CubT4vTznDZx7PTNah6G3o1PDA8gbU
n5agUuYOvUoQh+xPYIjI/+uK3k30hhIzxik4+wTuHhklOFGdZW8PrlxBJSoS4aSKTCeL+SH+ksUO
8et2EdGTktFpnrFEMVkIhzPgQDgW1nevNaGmnCpBLof0tG627QJQYlKXjzILTAInCLKL33zqyeO/
CkG39ACSaIv+oGG6JlYGzwCkZowGvn0Fd+Gem3ugAYvRNVkXO2/RQR80H+m1ENDn2NBZrsgBa3Ms
ahThgKKzy9t06jNj0rF4gCsHiiffVyYTW5E2mxt2rJWptHf/CO0zOwXgwHpvmqjAW35wpDkQjOt/
kFEfujSeyFxGbG3H2FONXMeas9p4rmYuPlsP60bhIecUEo9oNADWNUp0Rs60Oq3sBph7MTxR4HQ0
0UKKmymSCvNd0wHH6aCWtKp0dixY2VqdENZaKaUoOg54FiIDrjTHaRpN8XzWmx6bMKiT+aN6vsgr
kqtda3pYnkCIAhZxqhhU4OM5DXEZT+G6luQZdsA3xU3ES4T7NY3j1GEgNaa3VCbsBUuIYQsDJM1K
y2QfMgo1mtOuyJoldHlsZ65g0Uu1NeIrnOu0yCctwzAs3oiPZv6pj7oXiRlBNrAPXxG1sLl8dCXo
R9/UfA8+SwaxVx+w2ODd+WNdoy+AVaxde7ktIzhj3ntXhVQk9YwaBtnWXEfbDodnT2rdmlzkSqAY
6Ei+V55qdvTyVOHOmy34MkRlFUIsf/+uzVMsIVgG7PAPdpmJMqE7oGcDxegqkrNzawQbYaHaNHFC
4JC8HXV+La0Tzj6XlNU6GCizMJt223Wp0OVA/nXcDEOIISUhI96TrLBkd4CcpIdeURcRIjIlLAnI
j4tkDXUaD887btAbuaek49vxC4dAWWWwwpG76ciJJ/AO8TviaUR32Usvw4zGWFJLtw+A620wLxC5
yjrFr8tWBqwG03asPN+nJ0EbF9tokBfovvMHBHRmE/4wv4zyXGl2pAF/2swV0XF673cfHWJDSFBe
IHW4LQvHqWIGt7/mkVaJapEeai3WAL3Hh3kWjNxw0kcoVIkfw3YWGiVnwH15N6a83+GilG7W3Bzt
FzESGj+3Vx41pOF8CouY3CYoHYe8L3e/KDF84mEwzLvbRIp0Vvi+BlsmfBYI0+6UW5iiw5v3Y09w
Es1GN7wJpQK7esBTooqCnQmUeqHvb8gZJ8ETyNOTRxzY8W2a8Bl7wVayTkqYL5QvWJAdszJH6HUM
DwmB/b6pPsmevGOa3qyaoJspb3AvlF4wuX1DLo/Y0KWE5/bA5j6Qr88wtqaiz4hyGSm7g6ClYB31
IWWT3NROVrexmFTt9LGCt8+cYN/DI9SI3plYpsmDTFSfg4+b6TwO3PsjWt0wCBio+kK2CT40qsre
kAETTQaqW5OyOtr1ba6cG1epHVc3dxA9lTnThwjANTIUwXhTaraYYhHGKb1TlOubbHFixa3lqwSG
OGCuZeDqC9YnuuH9FlyH0QCPRQ4GwhXIdWtwZT7QaVRb8ji+4dKwBYFKEf0NbvS+3AQtFaf+l6of
My8167Kym1gayGE3LM24o88LPvp90XuFBwvqAB0ChrZnV0RCX//PXfch5t2s/fjlCLJ4XoPEmhft
GAVlqbxHED5oftvymI19vIEcnwrRC5wQDlasrV6Li0JSkAU8TttPI3g9+J2BlTPOyEwx6JIGxymj
Nx1PuVihDsCFDlcThfbXm+I+ahAVkZptyFEPCozM1o8B7U/NLwLTdLX12IKsvI9F4mWjT+IHBGhs
TCAZqnDsOGxasBr4+hux2wRGpLFwN0yDS/QCEG74D9CfTW3SIFRt+EdHVGRDnRQLhwiJsxZkxQ6Q
kalPWlX+vzwawqn+PcqFXO/gs6li3VVBOokBF6Z8+bPsaJzq5SVUs4s837+SoPLg91OVv4o9bpL7
tx/rEllC1hiPWohHC9EYWF+6mOA7mp+53lcK7g4jI9Nbx5M00faFJq4H0i2rZPACN77sMkKQmu2P
TdhbV4mInUodbyHv0vXNLy430ATN2LxebSDMS2GOjhV9ZvieWEbMyvW4pT2oEJManaxEY7Vr0G1E
0m2KzeUY9mvDRwe2uZr19rS4l8h2E/5qbcdLJNdIE+flhzNv2qyID+pCWNNJXcT5Eo1yEas/7ZJI
VdNJNy7OcEBfV+rMSqGbkoC1Kd9BCIn60A1pR1+J4jkDZT5gSaD1p6YwZdR/Ba16fYAOupILKADD
eVU0j0ay4LsPdAYP9E5Db8XmYKPggFJsKEvxD5Td3xQZqh3kC8KDMuhsyNwIsmg9nFH+hQ4PNZWu
PD1Eg7N+4tP5zlg+QdMLxv10ue74xSNtydkLcMDgDIHhyxyg3jahjngLYCdT7E0fabaslzEt0TZ+
TpZ4QieK06j9aq6b+IEf7KL8OBJKzniet+ZRTQ4rl9L0hAEvpfdxMfcRAX14WlFmjxWqQRbQWx77
2SWDoCRT1QD/misHTj9olL6ibaDUMtuz91FVQ/xAD1mOccyTdqnDWgMS2biSLHF3rKjRPEzqGgLb
hP0ArTO7WhHMoX7IWHaLBPzM2qXacExrpfYHcci/90qx+UTXua7M/xV0W1IEu9rUWsT50fBnIuUz
Z9xnwTWQkwCeG97jCdmlGkJ8BHaZZTFysFvh2g0rkIX1PBmHMJBr7zyYVQoMiY4ry7DCJ4yc4RXY
j4/qOQMNirz9UrPKfs9s4qsvxh//PJtcSwS+UBXAchuJ5O93OuO8U2qN4Rwhclc49mK0AM2eU0c2
M1twz+Y7hYgyvVV4XSvW3862iLO7KZcgM9+xKOXc9vxvRcu2Y168KHEYkIDJWXQU8b66PoVc4xY0
BenkiSnGUHJhsjaNB+3fzQN7mRdKcEPFnmEPrW/tKKRkG/NCO6q34O3zvEJVfb1vx40jsXMGYISv
6COgIkr0KX4O+0llWyEjtRokPbZ+6u43++UrmIZm0s19szusHgGeh5Cyzjw7IYLkiqAtV/9RkLgt
IYWJqh3g/zAGZmqtwgql4ZJ/PJISydBqSV/4VEIehTmWkdoxzPvQq9WvNZindmX1NGHDJziqT+ZE
jMfuHGSAB6TfIzEmL//la8cLe32vUfGHHXTPxGeOo5vyMjg+C+heGOMzRL79FoH7NjfL7+HNkK2Q
5x2gCqq/WcKK82dnTe2vKjeUDbl37iLhg5t7zuLo1W+r7eufJ8nkEaGv4h9/YwYYPRuMO+3kkHhd
FsmLqDE1KDjwY4L0T4qZOnOxyl2B35tWnmUXzjS6OPZ6bZLefieeNQYH7JzbxmOgJTqA0EedQyZQ
N/BFS2xhcaJkqLM45ZoQOra1aKhb0cWfcKvW45x3uv3Ff8hwFK6i27dC6HnSevTBfOnL+ovzFIBM
uEIowCWtJlmUW51GLbduEz+8KhicOK7G9i0CpFjemao4JkoMv8a4HnPQ/1OagXeqcNfryPKLc5Eo
jw+uS7LFlzu5wu4sSQXjozaPRfdPrb0PfIGaWZjcjGwVF1Lq4RMI8GnuES95I7+EgTbFTbpq97ho
WjPjZGbS6QGXdGl5GjOVTRXULRY2M/vO0SISu35mebBbt+88IZE59McFvBpCr8gHugPBqr/zrtFC
WhJCX1/QQt72vDH2jij65063Vu1uUZwM27iQfr14UW6RLOpsb58jpPAw2JKzHiCCeoajsjGZ6tik
5veOtzk95orVrr+2mI78vTaiXCJKEH4gg+tp9x9ta+LDwykT5fG+RY0CMryJ126OUJXp9yRrMvKP
mNrvp6k0LUdOROA2yuG/8RBwMkszc7TNky0FlIn0IJdsmDfrp4wkxfCcOzPcLDQhXGN3U6jbI515
DEDDyc7g9fsZqroB5hIotnuT9FQHzWi/x63hIYdoLa2/ZOL0iJnWL/YCDTBqsZ35A8guq/J8a8a6
OHpInlMC6O+vnYP+T64YVDrPoDodY/1fqE6CHsXKfY4tU+GnbomC0BgsQT/kc6DsUP3S4y55lBc1
HdeJdyaR/E+y0l8cqQ47xVDlWKmU/t2oTnrGPL908aU3agI8FipzFeEsjHRtJ5g/Cl3yNGsOvVPp
s+siuCK/WP7A2mPXy90lkcS/eAvjResi7aKn4Su8lglyO32B3+wiXRyeyFh6BNowHDvNy3ny+/1/
uidGYTaBqzUdyRX5xLpdcomkJAmL/Ky5qcvxsQsFxI8tEQOgS3Xzu2jadZP7yfyl+QAbJ/xFt0wk
5fIjZ/6jI/BlT+7iTfMgym7Q/BiDEgiGw3r7UEhNaXJV72CxBu1dIjXL7KQCJP53Mp8ZwTyNSfR3
WWYRFjUc+gBX/G3nIDcdpUo5OSwBXZmrgN/yzorOBCpx79m66Nxlc8LUrzc2D3pvpJvwxzf/zQkk
a7RxStiQzcpTWbsTBBEbF41T6gBgRlJ67ZISps7kkBT7QvZUP+xOxVQQmV/ZNxL5BBLcvyDzZH/B
HNqdsQ7WHhUQsYqHtBROgVsNNynXJVVqakhNRa2BkQXP/ZEp7JWasa9Jr7lrIxjIl+u296Es3Rut
p6k+XetHGkRAoXmOL0jz0U/W5V1vnCDIdTNmZ345y1iH75G0EtOKRciKecTV+5jzWc5AOcedMRiR
/jLshm/98lqJVl0BGq9sQNqezlIKxa0H1FbULk4y+IaKSp5dF6qRQotk8GCL6DymIoT9naPLXeE8
XdnANNN3AHXzP784zJIh7JCckqPhopJ7rmdpMllWAwIEryPNLgNwiCYx1ZjuIv3eNIFZ67H5ZlWZ
MXsaZ2LphvMIzT4Mek4EckSKfW0TdbTvgr026AlZmjP0jODyyYUAQRq+rzwWwC27XwJdDMctCgEV
vzbeFRjJNz8Mb1zgo4xB91rUtCDr3qYsS+xTWWBHL0Qmjf5z1tWvzkWuMe4dgmXt2/r2Bs9Idonl
+v7rJpVYNqomk8iVPtXXukKwgHCKU6KKf7+nwetNfGu/NTWokcZGnhRK4wNIXT2nu4xOphAgIlxM
45rhPmm1vj/q2Z8ap0sZDURPkg8aYryVXNvwUmBUe8nXjz3NDuUVaHKYUwe8wJIWYqCpxrYmogWF
UbAYOD0UZXSoFV1Dkr0DgTS+z1ZVnCLYmz9CtALmTqfvIxZPE+V1/8leWT4sQs5JxbEggVPXkvAq
XCcif7Ts1k1+sEIj5yRtJbDdRUNRsTTYCZnNI9gd58BjxeXUpq7SSlqUO22Qo5kAd7GLP8KlZQur
YsMDthqZ6oIA7miC6KWaWzhTBkl6/Ak5BvRhUxUKfGLGvsjcH+oqKyP1MBpuQncCpI0qtMCjRtgT
EOffd6tjkiuhiNMy3SRs7JKift0auDwuqTqoAXpJ/TBP+/VY+5xUgFufFKM/B6Z2Lh5HkT53ykQL
aJ0a9y32dNH2FJHURKyjekV07w2qScLcF2jkt3pbtt79VsaRbGj0S6QhkYhL3e5/BRBu99v0pb8a
EB3xdN1LZbY2qhBM0iVabcpDY8PvlaJC9BjDsmXT5NOFj6l3ZKEitlhDinAmTzVH/dCBW6sCUmWa
JtuLu9zyA//8D7KGWXxhGWvcWV4WplFrLJEMbd338BaPX42iTewlhnvQQdw7HbnXf/exsSFM3giU
pXj7Txm3tiJ9T6oLtB6IxudwO8gj6eu7wROogQsYr0tAAA88S+lYVcPCnA4IVOsS3N3ZeYlQs5/9
prbAt4ulaBE0zbtsX1N/s/J6WsSq9l+mFFXMZvgsSWB8/kAggEL9rwbeH9HCiVo18eX/CMy07NV4
y0EaGxw7V50t20loTSDmwnLQAL0NAivFA2raEfujcgloE9cS5gHGSdEUR/9971MCNyO1xLYo6V9H
eEGO+8C3vJYlQZgYEKEGQ8jGyR6nd8Ss93jY8j14v7vqeKDFNv29x6qM1brS0sRAYbZFPonD+rpH
aXXalCDN7AGvIgne3C9WJiu+ArjvNfYd7zvBcZAYWNTgpBmsjQfEZ3FHrwrcWdkwnQv4iTaHoQql
1MkNRLsqVj0corwo9YGGthIkjrQlFB5nFlC+loOQFFUKb2nboP92ke1ZPAN4UTxt4xVIB06rMTqT
fs093huhDbMsVqtCWGudYby2GemadRsCZaxoC2hVBizL8cKtA/O+MeqWzBvKsbYarVLjXT1W07dc
dGIXeFrN29rnYv7PYCARcJIviRE1kZg/WykRXKuwfM3BytQcvVQrcRmn5VqnIGqtEKlqZXkPuaAJ
qkQfosicR1crv2unA+Y0sAvgTneHm1eeuoX7kVDDd9rWcrOMqjnFRWeTmyymeUO6dEIbPWKoCITF
04ZDl9uf3GfRzwVpDMLFqNj1dwbX+SZqq1f4iacNQlBc62f7p2EtAaVcvzTxoodBj+nz2jbovi8m
egehyI+o5k6S3xUlxfXFp3jDpoBJR9yb38rnYBAhMMiZQ9HMa/mfd6z0v+9OainkmhQMjv6VMfhQ
aZN6tfbPd4vF4A2hN25hHMxeCBMApAGU6yGkKCMzkv0VJ8Ht2KvEt1pX1ozuJOv6xT3cnF3Twsi5
7MEF3dCPNXWn9oIklnzwGFx5vfaLYtr8hMA63CfFtlzWlBsH/vrZE4MMjSj/PGWBb08COf7WsZno
ZQnT8HHelMzUfzsWts2v3EzBtZUo5cEjtf9+3ANxmfk0IrnlF67QBfe5m6ZI5MbMfH4Arg/kN+ax
9yl2sM7mJe0vmG0g+xl6azYpTC9s7G35fIXe6XTdtbnewUrKqCfe2mY5OQFfqvembCqefFngFtw1
xnT+nJENH2Ws1besXnU1eK+E1izST4sJR4NgYDsO5v8SuavAmQBOR6zm/GDyLo+77tMQHVujmyO1
+wuCr1xg1hXQ7p+fniZuLHuW5a3wG5877NkgIsgEBCLZn/H5olL2GaRwyaV5vrHzX7d7BD57Wryp
nAC3FYakMzeKi8sPgXw98HwAvloh3YRo0TMEcE0Uc4IfnXjNuxbVR8rMg3WRILFlg53V1/ATuP22
D/P0l1rLnu3x3UfgbUeHCU7mrkjuVQtZ9CO2+kZdL4EYCrNs7esVuEFs4EexhM2B1K9Am5tGpgto
YvQkr38vWKVYnzNVvyrdlC+/YccpoiP3MRIQEXhIWCDomefNglDvOTC1Jqtu7YQHvAR4ssOZ2vv9
hivfXIJwqFOsmwW1YV/NRxtSJ2d2rmpkorL3kwFkxyMyGUutZvYB4ZzZkhIvLWa14F67TyWSZ6Iv
nEpfaETTMu15gOAz2IO1WDOXkADtnMTg3LStW7Dgt3MtWNZtej/0DCI8P2GPmxgSP/wQPNaxkrYf
OahrBk6Gx5rDWlNh+9JPgoHIHG890EvQu2mO7TuRxTsRdA1bgYJbu0ihQSNrCXliOlFKMvLenS/C
xmdit+gJ53LAo7XIJJmhjGgI1c/OB03RMQHruBnhEgnaaLIYZPEDemTZFRywSOn/AxvwZry+Po7u
+uWrHmZWUaI3xxZ0ILuTBKa+mAxzynLH6b0awVF13LtnmhY1T7clA7bcUf11162uMTjb8E51oA9c
aSQWU/cSMm7uQaTRW3PWYTgcQszy8AJVuM7cS06Egv+Y2s+pl8G78C0BC/VnYwKeA7O+o7q9tqdU
VpNhE0Z5oW2zZ1G7952BD4fJ1DzR/2/umWnCE3hBcPfc8qxkXRDiee3LMRo4M3Pn44Dy93GbbGov
y1rmstgxxyKDGRhJfDdpdufHWqTuedoJwmPZcj/cwJ//jUWB4EJVeeNE+k1dOF7bad39eHvF8UEU
9zYPkNs+lOh+SjiWiBNawPJ7R/KyezUpEx3DixqloaMtd7FJ/Ym73GRnLgOR9Uht5S55uQS0T9xN
woV6NGKF4fhNxlsLYsr9Gv7I1immGPI2JDnLB3QXlZz9m5Q22KM2N4T0Y0lg6Rv/Wi1CQq3jF4qP
mKCHSLneJD//2GV61vtgEFPxn0S/rohPDWtM/UHqZIX7pqyLFwBlqyX9KS2OmzXgCukpnfHKy0Fs
TTe7HnGmziuHvqpfb0rzW2/ufvXLgzpp9ngUa6R/J5+1yUfKNbp+IZpx2CR0Y9rzAfpYiah043oE
rWfseoSEgfDCy9ouIwT7VvsyTSos0SbENws3zJIllcTkByrlj4XIWKNRE9Ed4PBYhm7rpDrBrTp3
LW4LGkc2UZ1tvmEGnIugrjL87/OS2B1SvNWYrPgPqvesnl9XFAK6MOVx8dhb9kzMsprLoCtgOKVs
+t5kfyMGbXqajGUFGOXknXrtcIjbwrT1h+tWsPekZndf7LlZTXJnRYY5J9XwGFDFyCYy/dUCL0DE
q8jp3Xvcgf/HXIgR5W7NArT53e8ph2f7lVsxzcYPVt7jkPNj1pXwaaWP1opf/MjbQgvcZf42bLvk
U5F9Dmwkdln8DReVOCGjuHwzVqqlTfKzWcpEKARmC0W5lYRZlNbaJlLwoXpG3WFTfEY0dNbUYhIH
TwpWkvqy81JUhFBZjIs/ryS3WXG0Ps5lxsKq/jaV7gc6FxsC4BFjwJRHH9XinSZqPqt3ArxZUpf7
kYfQNzwc3bS/VTLief19tODlgQ3a4243BgNsXQIevUDDCm3xsXyi4n8oJ2zFkgpeAxcymBvpPO27
GnTcdqwcPhS0kdISCy4aOuE0iwFSAq1apW0xTyBdk8gETweZ1BR7Y7LsdH/iSfIWqKkHukgYRbAt
yQru/0612i1Vgh7wkGbshWSkNBE+VzeD2dzrYJ9lH3fRav0e5cjmVyMpiz1zblusR5Ej6aIIgIw6
XFs5OmkJcAQX98cPY1/DlFRvhAyhEuRP4nyOuR07+CA9o66ckl/qzAeTpPsw7tJt3TESmxU0tREf
8s58h3V4Ex9RJZBiM4lzlNpOvfxYGB97YBnpMvSKVyM+Ym/uuKjDUkG9Zn+/QVI5HWtYnaxenjaA
+anEby95segq6ymN9LRxZrifiGLq5M+L6D10MfYEk2yvZgzmWwOgMzwVVKHO/Lh1Sn2REnEagYpJ
YFvx+zm9EBpcZsE6JH4N8BvNUSraRkax7JNrhNZqp8EYkqnVayBhFHy0UXPmgwWfaa3VQ5sCnBKM
67svrPiAmKaKyFazM04AHTJn5obAFnyonZ5fYM1d8Q54+S2vZYdq3RU2ZWj0CNWOpv+IwfWMnddL
zsR3kmrCzLFneGhHWm107qZxmqNChsPPdiyhoKJLzzqNYKmvrFltM8HxYh9Y6fngK5DOj/en7/+S
h6SoMQmFywV/RH9f7wXLslclKbLdq9N/lsvESNEf4+t7TvJ0jAu3bCD7ZSGFuBXbEo4uFFc947hZ
6U0bIif1eHdfZ3VR+sYTCDjeORrYgYneLeqvzofWSGcnPgm42mz9lNXOrf+NRyVr4NXiCq4NHnfG
FXyM0tkhs5SJvGzxW4DvMBXlLaaU2+dKF8kuvj5Tx1UliUm3569RokGxmmTpiDjFBN/vecwiJe0L
zmK76uTfd5uSAk3VI9f/5rLRH3X2Q8U60HXV56FEOLoP6EsOSAset9Kb2adSIJX/wOTNlXnXPvnu
s5Ki4iglnGcqtZry+kILjjN1KgZHXOzH3wTwMqq3QWrafbNeXzdI/qlQc5MGc1nH+IUAKCxLJAn5
XnkHOxy41p8nmAExavCDtVhC/ry5rsTS1ngrbxoSbEp83jSTF4EalgaXDWetu/dAJE7bshN5VfnJ
3Kp3CeihBsU26zYCivNCGRSxJ43QpAXlaLiRyU4cVhQrbSX8+hVdJYsq08Q0Hxx/dLs23YWrOw/+
HqSrnDGpWLetlbJgz5nOOIuqFlE20LR4ITU57/hjmki7u+t+3O13j5A1IqeijT5g9i39DsZq8/n2
ReUJHdUsIc6HCzBBuRVXvTvQVoNC5sxbHAwqFXPSUEZJwZ9JsBv63zkxMfnSmEqFMlr2KsG3LM/j
492kxFhYiKuRUGmvl4GkL0yKi/Szh/YWtJx47Et06OOHURiw9JlEn/RIgVP/OpvyoOdxDCfLL6/J
vtNkwy4SoQly35vznAjGrC2bT7zt+lWQIhmS9/36PkL3VcHW5VH45fdlX19hd+MksrFnz4euZM6W
MFTuwQ71O4ztCNc6R6XPdN6cvLLY5mIDx8PpX5ILfQg3Sk4UmWS9VDeYGivAOasNXMmrkKeD/NNC
bfX32GOzEWm8iL26mIeAHL4XI6m1woXM573LPBjq2afpGNtG0UjusATyRgW/oeBhNyJELs4ec0OV
yRqbVvckwgDrMUM9pzW1T0hBvFg0nA22gKsh3QWTMZgbcBxR0fAFvanFTDmoE1D1WwncT8hpE+tn
AKbpYZb2+NRJV3vnzwzVo8kPxuvvq4XVq4Nx8Pv4h+EVEeKomjVDeeNx0z4OBnkwN2frNEKavYDz
wneLpkxpJD0cJ8KSUIqN9/YFgAu0QGBJ1c3cQHFDOsIbYuDaR7oeolt5FPXJxIanq9hhgSnRO4Sa
2PEMx7PVlBdVeJnY9Z2Bj6bTafcrmtiIdvFjLvRyiQww/8PxvvpJX3AKo2IIrrApbU1fevylo118
05AFczLdExqy/CJilSGP7g9HhA30Gs24hu5zXPgnOQQgHGEg/jcI9kXvu6UAGETmMZg8dkvRhi8q
qTSy66ITwQczK0JdRyyLmvGcod7oTdIsyO/L/vqD0fyzwLANvYkAI0PAgG8mMPs0fQWfblOo4Cvx
UuHdqTG5XTfdG9USUv54kZrvOURUDwYFwC/BHe0gHexdQO3tM9B4OeqT0Fp+qDio8kZ3bcdDrPPY
4a/7zE9gOnAwnrVw+W5TMv1DgFPqKobXfV/2Hiod2YNe/wnZcb3KxbXXeSnY/k3+GBCfBPGgCdSD
JBFX8Kb2oVFVJY4pmyM9mllcgFyVUwebFsXNXPBWmzrRXoDMGoZz5fAm3E/VG1VZ4CH3qHG04y2V
G31pt7+yN5D6K4/4bHdBeMh7HqKqB0c2yNISIpeO6Jl/hJzQuEzhuHIfkjt4pZwBWmf8DN8ofjLI
lYmjpWSTW/woNxEAAMi0L0NHgBBC2i51SUuK+ezi/1pdccRg/DFjueOb1wimYeS6qknNtJYIBuy9
m4Bm/Rk6t/V+gnmOGC0tog3orgd/kcOfbb2izLz4M22S9JN2jtUZqZsWvfcuKBvj8mIx18u2NuFG
3HxMcAejpLbzqNKQD0WJALFtG/C5hTWutcznLV2IAX1GmeWsipoSNycQ1o1lEXVBYPzObbRvCyCz
tXMMjO2fdGvPsRy9p+ubeHpHZ2Kh8Wk/VuWeCcYNKTiSdytyuxBK8RiGfUDp+4uSGWq0kUYLM9gr
l+7C/jIAa1YLA/cpa14drFxfBfZDO1WcAvV/21zG1e2/tIGl4eYuFdkb5j6q6L0RpbpdnP8w8v/X
WXwXqkT0DYpV2/rLv1l6TwbknuiWbwtWOowGzjzkh2v/1EWmvXKyFIn5KF5ykdnj2Ho6ptwB4zXX
Il83kDiMUDG42BxYFzBfyklEm4nJ9WKjsqOlOEBQC1o8/bNdjHtKZW8VUgb4WxYZ2//S72lQ/aR8
RfoSqQvD7BdGj+ZqQboisulhDBPRxY2LHNselgYsrZYSjgQ2sVhheQlSHBpYo/92RuQKVemLN5Ne
MP2vsv+tqOraYRMJERT48rrGXDdUZoCFob+/vArN0IVTC8LMvCttn/uCGx2ycnf0fpLu1IkmEpGQ
G++97r9R7rjzyMddpyJrftcyfU0t6Tvo/OF6g53j3WykI4CIbWIBzlHOjFrfo99ehKD6FAshT2yc
Sk9w2s/AZSr164KRUYSM1t2yNHPdh/SPVj1uVvB1NUO2y2U8aWY0bpPvIi0/SQfjRY6Lo03FeQvO
jAbtD/Md1U+yf3VoHWugFW/2ad/bEvPk4VyX/V0hxJ11wzIxJWFoSYrh7TAUI+r342sm2/A+ytpv
Q36BCAj1P+Gncu1sxlZ9qLANzohHvKwYPFbrBru385bqHCUhzd9BkXWu7uP4j9ioW+HkiiJkcZB1
rxEhA+XesRYXx4UVabBKT2PLv5/aJFBSJl94V06LDOGuVkl4AY7OOaDPI36NiAOApaAwX5UQhZ0V
9fQr3LEu4h76JaJ0KyXvqtfG2+Pe5uxE/ai+vfIPokcs+Wj5BK6hK6b6gvJBCTPCsY2GjXCZ5NyS
IX6xSfO4c9Y4Vj0gfx6VIxpQ/AYduoEFhtzwGUyacBcsYIl3ZlqGt3FyEOYhaXV9Bp19o6UKyy1K
/eqRRZVyzzE2fNffVny77PsOCpxGDck4JtOuswwZObeU8p9EMXY0xznHOyF0y6hLsneK++1jb8s7
5G5gC/YysGZo3hIygKLCJNz0/Y5e0rbROajgc732hMtaBpEedu8L3R6X5ARor1R/MlOlLIxZ0zFX
9EHg5T92GVsp5dnBizCaxuGSE8Av3jD59iFugLi1cJZzT7UI8ufJSdVgKlSDeWp8LpleFZ07ESjd
jd2C3j6FTRTvzJS9aIh4UUuQKHcy5hTZesni46UIY+1aP3b5djOdC7KawhrN0h2ifBlRnEXX5HPI
clCtheMjR2YMlZw9y7Me9IXOSXzFzAwKa87zEc4b5QA6KTDaELDEHumpoHcHBXNGEJJTDV6f3j5Q
VU0kT1+49FvhDMmFJ+6Zf7X2zNE4h7wdg845/piGG8pZPeWiKZQThYMh6H18XWLnfSXFxnsv7tdm
Zkti6lyLSKs8GN2YxQOlhcY3qOWSp/e5ovySNNRi5hdhLo93+4U4Vngpj3vux0bVHriSvh1Uf4hZ
0lQWwBWnQoRwS0cRGYL3LxAj6G/kGiTq4v607tFgbypiQmw68oZlMY7yyqFB2FpbiK/Xxm4jYLyv
wvHAdyibWcYz6EYnDUhDb9dxYr7293X4Mfj8q/SN50/aAZTNZE3YMjAuSIDuRWNX4INChgFuUIcr
64/3P1bCdXGrjOK0cpKq9dJx+PnwmoFrVqWR9e0kkrD9whd+1inDfuVDnACavKueEpkbcEvHnHtD
3vvc8rpYl4jVvFKOXTciS0eAYGMaGVSkesqcyPUybUPSzlHbYc0Mlx86K8Dq6UuJATHCem5UraNG
o4BXRtM3XFciutAnNNkp07gC0izRP5L+f1ZtsDNS8EEuVXGxoV3FTRJZDxY7pIMIgmEPzRmICyNL
X788W2nyEFhClRUeyvHZplXs/nZVtnDFYOswDY4joI6Zrj53Wy0VDGj+Rsi22cAztlEBdtWXbyoC
0Txj7FagjwWXI4H0szHMxnYAAc/vsDIkycS8qXzBlVLhd9uUwC1Tc/QQKkoiLRYgbYMY7JGuMLrN
GPc+ELeZqWGxZD1rLzqCN3EIiL050dGmOBB0h2FSSZSL2dNwNDBVqZ7/IBLmbwbGUcq1qacFUNXf
/DN/G6BRk3+QRqrEQwnGbtLM1JeLpCNRfbMmlJ0YldfKj1Sod1BZIKIGKjf+1wCb2cg5Zb4TQgQD
Di+y5ODAyPDkekT/Ks3vpsUXtPUltuJf5GhUUhlP3+L3+RXZeON0LAMdp/CoFARFUlNTMN3mov7T
eed23gZULkjXTBK3QzaisVSAzJSjVM6HEm7MyfKpeGj5HBLR6+n4T2IM1pqjydD0xvYzzHznkBQW
JKGqUCh649tpYuAIoWUkbya3AfMVfOe4TrBbNnsQL98RThpEjlWxySNBNH4lb/OgbNcPH+MhS6AP
8ByvivpF80CrOS45b9wfoz5ih7QVQbW5LZovy+n/oB+KkbMOK4roD0DQqItC5K+xyQjfUbSSzzV1
CqrEGK6ch9nOWKAxsDf3RNeQsw7YrM2uRO4XIoXs77L+ZGN1H+TnGCNFbmcn9MUMi48QlT002RYh
NoE0BiNTAz1Xxx+a56nqEEbFRwHkdCK8FhAxbYKjfdlnj3LhipoYQqrpPLpcw5GKL4Or1fPb/9ud
j4MrRa1iFP1GO6qtT2lb5Q4/f6ESKD/89YQagfNqqkkbc5SKPV4n+7jJLuJSeM2gLFp2uV7NayCz
868J5nCiQChHIEOX8z7zDjeKPVkfoj5QBAKcR1yExZawWjegSYPHXV4eMnAt+vJbQny1T3GRDm9n
qb5spYnr0YpZS/f/4HlcSBZ4L1BtG5Mgwz6hb9Mf4Dp1N364ytg13Zh16wuxariKjWtWoZcRjM3B
YMpIH4wiKZiRf2K7/jUkeRydw8HPURSR6Oi6ZSMVzR2QZT8WZ9b4kKSFQpI29AxqeudlUUiBcbU9
BZqcmvDeOZGD27Si2ipHc+tBm1i/vb1boIKNwHAtcx+KLxmHHwCPtuKHUizmFAauTpE8kt/rDjFE
G8zHQ7HiJ0an5B5zasVPyJFrfDl53sjoIAsJLr9diDkuexaTiZ4K+gB4i0/z9C2BwwdOfOi+80gm
p74MpUN8OL/RNeir+BYLktwOhXL7PMAHwBqNPpGEtg/yYntvlwcNEVQrNmuiz6/RAIlS3qRXO5ft
aP1TX1p6p9vOaVWQfy/ngyxFG3HSY2diuP9LV/ZwNw9DvMjAtBDBxEDGE+yXeczwQ6OeSJUylo0h
ZdfOA4d1OX756qxZQYi9hAsEoz0+txi70zlJIHOaB7x3RBGe519x5dDjBoKdPpZjuWTaX4ydCZ/1
QqHvVmycc5xh+/dMawuSISV3rx/o1SNNbEmknSi5QI9FID9ZUmLjvGtv6QesBioNBqQU8yRSj4/U
DGpVKcM+tXoRlqBWk4m0FDem/L5dq48QLXE4XcNp7DLpkFO+Jecg2FeI0T0Mmr8+bTMd37SRSSnY
cBdqmNI6BxreuRSvdfh/jvCnXq6dpQ76amSF+ctkCEg9Igb8SYMTnPcmhiXlfCPd2nbbSqlWTuo0
r0kD4SF5hm/9a3Uo4tlocOc2rTqJOsp0mMAUEWUj/11goc5U6npXAlkfa+4n/7I/stgr/lgQXSYC
bNQUUZQ4ZkM/EY3bnepoLc2E1lN26eGBuqdLsSjF0QDqdWkvS+oz42eyeFRthX6J7sCi+TFhVg4R
WI5W+yRHWGAsEQBbHtcvEIF3btjhlR6qWDCo3/4RXqmyPcmPa8vhooUmoiGvaqMAXPixfna+V4Il
60YK+b46+coivlxQq4ckXQr8viZkhgO7ZK2bkgKzO005G8khhFQ55Nw0lVx3RfvYq52fNaqWd/vj
QxKK5g4oUNaeSsEhw6W56LblRiQKIHyyZ690fYVHF1D5tvdo7KZw/nRQEz3HZ1B++oFOXfefLlx1
cbRAEbW0yECb4GMYlVqPD+t8iN/kOPygP+ZaRihzeOJPiL/A9YYHiCti50vjft8NFOzta/F/QIB8
CQc8whacjG74enxOTSP0+eA5/eVMLzOZXsmRu8eUSkCJ2WEfbSjt8GqnkKN3CVYPDs3t9dXaa4eU
ZNab78FyJP/zMs4tCYstDOXGyEdohJPmszidNnRscAChKeDZylnv7JJ+cArecrphzPczSYhURBrT
98BBxoOLL/8Jf7rqfnv11DUd2PKD6EcEFTe657Hl9y4Alq0ozI6cY/1U9gQEQ0lo+ZXbqBzm6wGa
RcSYqCeIrBkNF7pQH74AEK0BXJmdZk4T0eZtG0tSg01V9gpdYTngKOfNeQzbxud0KfqYvdWlGeXT
A8eWc3Wlu+QsrLe8CoPmP2odDZk7BZ/hwDgFPTHvU+L1JeIHtEg/THo2BLeIjgnsoCPXRlQhivj5
XVcabSv3lLs+WpFDqhrEa7JhUmfVTaMYJ33GxojLevvkubaX0k5uTEopPmeRxDfw1Ruyh8apchfQ
1PG+MTlQ1MQmUqmHOZuhZJOn5OO00zk1PajTFaFC8kii5wYE+qVfL5IsEwtaliFqrOdo6rFht/SS
XuteEF1Gw97JbG8cZypN9jN4zTAUnRad4Fh6hDV/GJQLIhnEIWFrdqO3r8Urew+5WyuOs2Mf5lof
A2xmW7ZKQt8Ln0SNzGe6DE0A0ndVHQd9swUARzhsMuQ4/x8gH37hKIE8i0qAlw2ixctaero5Wiul
ZppWa0vxJ5wwM4OM7mFrj4/1sCMkzrigiV/E9wX9aM9GgQouYHLdMqTXU32tkRNoa+16uQ9A+YVE
cbcIamu0qW/de7OZlmBqQa5GU8piSTUTTVz3eRfKXeVdR87zVKyKh3RKx0V9RgCvtElqHC3iKOwa
I1zwbtss2fpoGR7zonVxZ58UWGe3oXlTH/q/HUWdCM435dJKv+tHgW5DIRz/ofODd8ByKdDxIJ38
xiyui/tzlSFc/Lgd2k6DXWp+WAOTZ9FpiVaNt0hZBfUm9DjgC8hJZSwMZ8aw6TPN4Z3a6hX1dqsj
DNA7OFNEURy5snB788TzTsxYGbwX3Z6pQ4l8dWqU1/L0TwfX6XmXRS1ygKIjeOyiFxq8800Yeke6
vqC1MLxUQDCUO9mhCK9WVAsUg3jmeoUdWILtPMp0gniV3JfKxXlOW3nk4YP9p0GnBeJnPVWAa9jr
uS+5COcDknU3rB0dZQXoFCRoNv6RV+TPiRTurFBo8k6jzIaaOjmauadnPA7izxwiuzVHDN95eqo0
J6iiN0/M6XrvGa05I0KpbXR7mohni4/J7B89z57q7uWzZetuVh6ipBjxgSHUdzczWzRPiOqM6+ga
shoSXg5TIpWmVyIP9/ghEXHBuiTEndKiZM7teiQhkbpOreuqxSfjrkpSOgmRBTWkBCChQBiR+QtB
a0od8AG9gqXd5r12sHPpb35Ln5IyADF+GUcNM46C0UKiFKW+lmzyoabiy35sNR1kYSxeCMaAepaB
i3a0cZfhmn8UyZQr616VGfdTNk9FEPf8l+MhOj8/fo416nirZbh4A78rwBDyrHJablxMrUkBY7Ps
YKr+PIyTn+Jb1MuP2hISvWGXEuUw35DgZzqEPt8CktmwaTE5PZIdAIW6bi/NMPRn9NhTKOBc7lHG
Be45fly5qZhM+xZlICQvVtGZfKtb1Iugb/95LZMyT0foMg5od7EgCeBaCHMZsv2cW2bz7bE9i6rN
gBIEpe9/KZl62P2vSkNrYSiOeaYDeocuy71CGuQtCCqAh+DLVHfLGGnht9Z5n0bXn3gRZgUifUrb
k4byyHcLWT41HReG3JnIlks4vmpwPjc+vulr2xOQ9WLoBXK4fDKZ3s9yHWu3X2MQ2YyCUSAM0H8Q
nm5Zr374uay9XDcOtesaHLhK6Jaj8h2cgLMmuDJP4CtRViER4c3ckI3h0pFsOJrhoUVLWvOeGJsq
Y5/9XnR20ztNqOxRTpWNrmKqqZVFbPQwf9gEzR4Fm5DLyYSe4mXgTXdZGASja9uijT7E+Bx3kg6w
Ulp3vK8PdSbW13Vn8oVOpj3YF5oXzSAQaLXu/JFAejdwMWFBfEJr0G8XMSiTXzC8QmXoqNTw3lpS
Bqh9bptsq5vg0xqVSYJeTEymEEdB6Tatm8C3D72K2bUtZQQT7ocrYgzu+xMGbaT06M3cQN0tWhCS
xUdbdkGz1YJdxc6RGVqlWHNppACGqxmKclMOHGEwzhax6cPcYrVx9ufAMixbSy/Puq5yd7gZykBO
0r+H3zIyMrsZxJ6mYyBfYI6YnLKjMyUDoeE3w2q0EQVIyUSrE8z0ly2qOnZQmHtLREKC3wGAnVA9
aBraxxf9H/iwMnhOhJRfcAmvntShwtD3GPUOcPzLDVYinGhHlfkbrK7SAtMDCqZgPS2QSUnwJ1DA
ZYY4QXwd0SkwQ3AP1o8T/VmlWmofKWepAVSXn27GiuOb5lvyVwsooLo1vN6jbw5uhcGu1Gqj9ui4
6oUi3rm/QpJjwQOKvkwvKj7el4ZSqnj7DrMP+bcExRgRppizV8rF9Lk7gJX8fy31CybvfXiLwwwt
r7Pe6HL9s3ujj+UBItT0AhYamL0stYAZBXIGQTkwohMZzN9ZkFLLQlci1HUxU+IwoUoo3KcUN58O
hLQU+Z69mzBoic6nSPxxbdPr2wFrUM5f4k/WJPStR+fP+Tn/u9jV73DjThyevv1Meft2fqeobOUO
47ZUGgiAyL57L8FmUCtYZN0kl4i+ClmR0qZT98NFFTDhOkgRRaSCVDF9NkWk7s/ibpVBjE1R7EOK
TQeiAr7CLHmregkgGMPHvFSm8HgHBYsXgvVIBHEf1kJP52WWpE/uQ5BUIEt0Cy0XcgGxBrgg3hvh
oyGfyM4B6RU785mQJcYbbu56/yZTCoz6vcMTH7wrZDTyDTBYs+6ZL1wqoLDc5JZ6Z8L2koPBf8Ad
YIVtJSq+dvVjjk1XH9UQHUyNRponegH24Bm2j7zRqETWK/KaCIAGoMI5RnN6SZtvF7zJhGrwtuUK
pHZ2vWLXNFYAHyQKwjoP5txvQpg3YzGvEtwg0IAxSnUSmQuKY/u5Xh96oAlskOXnu+SSHQgsQ+Vd
yovXE6y/Ism8rpHBBQCLP41ydZ15qXgPH3YIx9SM5EVyDkRlMYA1oW0jJqCmFi9fbNTp7AG2GQyu
jzRc9UrYkvfODyVtczJniGeez3pGm2qnt7Y3PxCdpbaz8VaFCk+iXYiOjEK+3zUUi/3v1Y8pZcOk
KI9I29we56j3JdVqIWQaYxLwBC1M30Rq+fxCwrh/RkB4ux6FXiKWy5MTI0C9DcUpmsBgcUpSvOen
r+lKhMRfWYdsSmtCkxgMIHZ65BHa6KcSxjdL3jwrRE2PUr4w2W7BdImZueHWbBzOuQCC/C9hFsMI
Cscc/gh/idHCXjAz838SWg7KT+sRg41upyUJEeghQSE+idrW3K/EDbk9SQxCrYaTl4yFpsPd/u63
mAXpK/ZiXboPmi2mEn9ZmNlG/uI6N/wC6J4On+bjZFkHYReMak6JRNJNvqhyVNqeHhRwi9VMkrrg
BFP1rhF6fpn0hM9IJns1pkUgLppSS7i44Z2ls404ikEfjBZKpbvTgVJ9H/8OmAB0Nc+OUuoF1d60
A2prjLIQHHW9IaRfIJcJUUNA5jk+p0Q36cMTQmPVhBIAWC7yUk2YvF0SacMrWmhi59W+Nm470oO1
Vga6UOeVVV+s4YLgwbqgiIYmlxVotNUF1oToFepJb1b+tjAnDGLX7Zo3LLEWL/UIVffRseZSkAWb
Ee4By6EdD0fCbTabsnu9iERzhDDGAswDAtVJLWARl9NJ4wvpR96OfWeD9SG9j+3y5/DtbcZLsoHb
J8qoTKgEsNCS3bVg3mQwTYfpDn4lFHx+djajDh1t/JNOd5XNlo44GWHXel7o+o+L7nUm4rJ+Z1RU
WSuCakqRdPvUHECyghFqEsMOOyRy9XaCEb+8+NK0Ymr7h7+DGbXzkSfAo14T1tJ4ZBSlRq/5y5NK
IwrbcxB8EW3Xc5npkfs+wLVuy9JFnFhYzSeD8Reu/FDo2hOThJBfz11enstUeslHFKjEOFiYX/Dy
1bnbNYcyBnyZTpdVOqxTcT77Zi48qC5J2wfGPMdRmiShZBX3Ul2ZRxuvW0fgPdK5dpv6rY0YvFG+
7ulog+Lz9XvYTog7sbH4DuTD6MpYr3FqT1OC7k8L2BOS9VBzaSHzlqzrVvydLU0xT4drvonmwQNx
r9t+CpDC3nMwTWwLTx9h0DWmtvA4lUXfjpRR24LPckgm5QrEzn1jIURFtxGShnM0DV+k0aFlikbs
2c7SS4puNEGoTr91QbiwfMnpl0tHyjn3BrD6cvckMb0ur1FSZ2BjlPmFDQFvZ7vUvwt4URCFnHCt
ZkD0RKIDJnRHrYCjl2b/Z3zic9BdtY5JZDInm8iRCKSzyYap/VLFU74PxXMu9EcWEtdwe9AWMHRM
UBJoH8p3hDbebb+IwygbDIwc1OhAotUzZOc/AIoQ5S/0Co7CbodARed41L49thk7HbJMY0HfPzem
n8TEQ8Fo6DTMRtEsx28tdbG2q41AiYjoD3Fw0b1ztNsC2PP5CfPD8LQyYnrYflpYiX52x96pPvbV
jDBKNebZv6xijJxrOVzUMGbJadp+EqLfSTuHjqnWQUKI5eCQXwgM0nOSVo9LRWMCTIt+/nUecYzJ
puW6IatxF60sG+qa1b+vTcB5BpTyq95BmHxJB1VTeb/YQcwH/Bx3GL6xRadOpMhvRpMyU2ZHsy9Q
e6p3vIHNY60ZJ01q7AZOE/VVBfC1cdgvvBTpgxw0JZk0JAg6f2VZC+Cou0KdT7FAz/Ng9oGAiEjc
xK9bkGRLf2wifU8S60rmX/VvgO8wpTHpKDbIvpu6xty3HWfqXQfb9KHDv7P0Q/GJg39J6K2qOqWa
Q39DysV3lXxE83WVIeCth0CD3a2ru4sqdgB+8rN3hCxFpRThOIEw6osMdN54rupfIC/RNg4VoOKY
qzIiBZTZEW8HcIewJQvhbTZ5HUpGGc1WL9Xwx8ltik6pNqm7zV0LuxTxvZEPHtZFNCOha1En7dbF
MSK1M/JHM0Nvhd0FV60FZC9YivTSF/E1VNQvyX9bTuGfzWdk5+MHa11UDTMacm+IoHjfDiVRmzB5
lvAIx7A8WIiPV6vK8CSKB1K8TlJLo8kpZvRkkry4DHQcSoojpV0WrV3zy/AKCTJMzZTM85IjjgnP
2wUCb6QcbcMzlnW5YKs1OEOhr239am5Fn916oZyflPD3pFGnpF8ZC+MtksMyYvmEuutgvWcdJ5ee
j4WdDfiVHw89PNdEwBOBJ0DzMXRpJsUfM/UFiKnrwUPzolGr9plo0bcg2q7j16Hq7yBpbwk/TxtW
IE+KtUEy29e4JrmVAh75nAp3dZPY3bGSliu3393y73/MvVWTS+quHowIFGE6OjLSjP0xhVI8pQ1k
jutH76aCuVYpf6skSw8VGsbzacqKMulyGIOccUF35W+hjgbJ1SqgEHphowFFp+mjyAdqeys0c4/q
BmuhggWzAG4ZU4Lat5/9tnHS4NkBOgix4Xc6s31ifKrAjBaOFyNAHYV1sQHXDwmqKyFrqlslCJcr
UYO+obhTXJDFL9kt6JqfR0eP0BUT3oB2RWWNjruVUZhd8vbUAxibVmvrqu2rT3M6LtdIJM0rHHL2
sO9ev5zsNHf0RCEine9/9+9EfRzXMvPwn83jEhzLQ4pGMEts7YMYXJSatUui5Y/5DAboubU3wJQs
4Grs1bXhLV8JJmwnBtauvOD8AU4yNn7jl8yvt3iYeTVk5pMbjKC3qeaolmfxTIdXBBoSXtGx8Q92
QYhbI4aHgU0Fj8SkOBS4VTpbSmKvhkMR5NOiI1ronFR3l4MQSt6PnR6ZpAPPxxFeysPeWkI7jTeY
CdiJ4n+hIsZN/yUK+5dguVVYWLdhX87PhVNQrJnU7+951PVEx2WMhhi6HkKY8SQXWyRAvaimeXg9
n3a4V9lp2J/zIZWAkjeHjOuujX688eb3+WTccw+/Bq3b74yCxcM/71jIby6IwYFa5Fb6BE50Y+sI
kmqRyWBKYJZXL4vtBkFqBIkge9Ce4a96a9lG3G0pu8cuo9SKoddXyCddfU6NarHD0n0vtY6Vo4NC
ssFjao8t0esZt3j/MoZs8gQ78fiUDcjpAwu2ChHJDmvm81vXfsnBHsQlSdxvSzPNzwSoDdHl/ESE
DnKuDl8REIuE9tLS1bxdXF3zHXwFBVmaBz7DB7qCa+0pNmE7xQE4xjkYDzMKDTW/3Oagrj8EgeK0
/r8pUXaRAOj1dWyUrETsI5rPoF7w9mXefoh4s9Z0WlvLoISzXZtLGutJAGhn51AINPYrSjAdqWWG
5WQ2xwQAsRxFmpr27z46Told1CZdKc2C4iiI5gBCQBjXLYsmDIg7s1eRv+eaUdW01IWRE+tITLud
Tl7ibAOG5rolA7Pc6vUIFp3qzHwHmHMz+2yy6AcQTQtVfaq2LJDU1YOzTY1JxWu0oz2HgG62PDL/
3bWKSwhIoGQRwIhTygCIwnWnOAUVY90JSpjQYfCFKr1LsPjqqYfTB4aF0tHarkVUB6/dUcuD836Q
faG5qtkKfvVgUvivdo7pbAHSDb55tSLxwcIDZ+iIDX6ITuBVYbBUrDlxrbSsBi/M2t6AHIGMwhPT
jy2BLFgPIbOILQ/z8rF1H7IRaV+gErSC2dPtUkq7ghXtqb/2FlOMUugzbUdc3exd0Roonc1QY5IK
jE3I5PoUp/MKqwt7xaM66odBDPkXfOxxVzKuK6scIegt1ABl9Grs75Rbzgouc5SQxbwUT2iKujgd
QUtwYLCkoPGBZP+ZqDhEPkm5TJAjsLrDvlgzzAT0AByHrXsVtqTPNiUgFcpRqVAKvXUtPamZQhrA
P2J2JSf0GjWKEIsL31y/x5j36WuU1/j0esI65HMmay3GeccnEL9GT2z8fKJNYShtEHpxHFtqpdzj
0zMFidtZhQMFpM+jZbcZqbTue4Ot0VDbs+W3JufjALfJn+aLFrQU9PbMRYHXCuhkFwiOn+Nc6B+I
9WY0mmo1s5ccSEvG5eOHX/fj8zuzw25bzrHt0zc62kMqOgx2xNN7v0/iNBiu0hBnJy7FXUH3TUe1
RG3fR9c1kOd+kdQuQl9QeGrAj0LfoSW6CytyvNl5xV9z9QBV6eekj9eA5038rzZWFS3vicEtH9bJ
rdirp2+bEusMi38ab42gf+iOkWzssO+W1VebY7lLiHhbySh8IhAJjuJKf8KFQSedxwQnAtNViDQF
We8Yn2Jgx23U60Ax5KasgTutuk5eTaqjVCxmnit5t++DlRHRpTa6uhDdG+9qf0+C+MEnZNor2tfX
PFS8wW7//elpgx6Mvlm8V0zur8tMfl1nXIRk6yMs2EWDJRy0qE7h+FBzBPPJyAjGY7pv6O+MgBpp
cnmxiMN+oz3rqnAkZ1BvhJtjr50DH7YUMlUTqE8S3w9Cq77fGxhRkIl209OuyKk71WIkrenlyJqF
1NxpjOMgDt7ODh5pTTUfeR2WBggUUhynmD1DgznroL40ZqKOXMkiI0W38jaNS6DYUSuL1Di9hYse
48q0Zvd+Z6bFg79EoYiBZvLcRkxlKz7UPWO4BS8WmGUGB7O2laqp21llwpp4t8LTAy0nq2SAjfrC
6iSMMVHawxFefpSJ2Syh7ldqgXURh2lRulx9uzw9uSjpGLik3WKVh7Dm3hir4ayyKndqlFeDjIxa
LshL8FzVKWdtRL4UyMVi4R67AHUpzrDbfv7AnaB/lfkGmKGJ6Z5RKlfPiA9zIxlQ+X7habmikK9x
ULrj+U6b87rQQVVHttC3M//AVX8AYyE4f2l1T+9TWU49lcZRpl1RJ0YPg9VD3foTrlYW6+B4swYZ
JTHh/CvDDe6strMYiYCAVCYtB8/IldZRf37hoIyMSQtEwl1B78FkkeIFRuMGT/20QtiL+aUAteYV
BUFtx/9mhfnd3SJU/GWhqQwDBFX5QjLBUMNmAI+3He3BR52Z/ctropUz6EEhFkZ/dno6c8VmVqUi
V2HUv5noVMbRkfCAUvUVs9iS1Mb/eRk95PFygaWaEZeNaSoTb5JpcEK5DQWlugdeXdjqLVdWthe7
bRJlMTQ+T8xTQ5Hi4/Sc8l+LlQr3YmvYRE/2ccMhbHx05GCXrOylzyoi71o44tn4K4W9E8X2IOI6
iwr901vUd8qrnjxXaTQVaz6svQpvlLXGebsbMZi36rOE16fV73ZMBmRrODHEEDdimil2D03z8dg2
TSbSaXw+GJJ/v+vxAeEd1FWcOxudM2igpKs41hvYvXlLm9RZZbmInnHSjyYD6VVXO9Wz0GBUmuM2
moNOqyX3UTOpDYzlg9vp51YGjmIZd8y8tl9uMNbohQjggYfxbzZJizUg+irRN3OEBbTDfGlUW1Gh
4SMQqzXXpIUk2JPrbjwOy7u++y7BqGeouiRZ/N/KsHcwIgL237vXviicmA2xEtdeVsjntE+IPbMy
Dnt5tgA6ZM8qUG+J6AfUakThQ9lxMT/YQisS33KX/PQTRtvC76uOT8X48uSV65tpMJRJj3J2h5OJ
bO71sVJsZRbMzpUblNqSgDWPDdXwkrePxKCSIkPlywSLX8TrE6CuwzfLtcusTeo6OKTPV6HqRtpC
mYk2NIpRxJlS/IWtOFOmpnNDLvFBQNK9CWhR8WCvr5CK29obVQEvV7S+DgewxXcFpHkRT2dpM+T9
8t8wH3ai/5oGKALujNhglVcjr+uUTBfu3IVx2m873lQlrOXQBzB4fP9VMwQxIn/IRY6s5fCs7Tug
3C1Py3oPnP+1rZdlNsPK89I4dZKmIyhI6664/cERK3An3qI4tb8d6SHNMrfQN6HTgVIlTVrVb2Ra
gEAPCGkaXS+rpc0LY4cvVLUuC93+WTXO0bdnXNGpWIo2q9N+eQxyFfrfEeQEgowkphblELaNT2Bx
fMiEG52qiDSG9o3i4Hii7ft9+EnwBSK3CQdMpoTNKwhtnYPU+cHPV82VDgBxsa5dy0OKnE2eb6YQ
xEmRotitYSzIbxAuwl5XKTrnAUTYwMcWpMlEZfKPvELAqonh5Cj3htJXiKoC/M71HepsXo+2lKGM
CPFZ0+Z3GypfjLfUl59UqsBC0sFhEA+LQA1Sg8u1/v0pbSY28Wqv50Xp4A0/2LVRVEZ3caEIYrMb
WSgUiZndD9JcGoLLjXgEgdZ948FZ4glj1GfliP97RBFqDe4fh4zr1FdhY8fiIGN0ouzoq5+9Nz5a
yJetW4Hx/dh+Q2SBdhpP2A3V1ZRQ+KdISYDuQYPMiXXzhZSMQ8QyDU0vx9HZ6he+RBf0JRzvQALp
HvclbP10ICZipDWrT+5RfsE251iTn+qsHuSEPqMbnG33a5rF9ESOEM/g7SttowNeTUYY/NyVUmWz
SO0gH+89lCgsc4oSm6Qvh7EXZGn3qTsNwcSBUgM2z8OvrpcyLLcfiWOOyn7WnbUQqN1cwqabTDwd
Zpi32Irkzq+iZ2Lw9qOOUG3yxCfQF717JDYXoMIuW2JZ0g+wuBPVJhKlpoTol3dEmn7prjqo5W7s
YuG/c/15e7Lo6sNbP1De54ykb6YwafNS4ppbdHEaJuNmlADurOJ2mczGiExi7SuZo2r2/xLBw8qh
ENz/PyKdgSsGDQIreq3GJ1/0yKrpNcbyYHpNnq/9lus36uCA8bINC7RAewAWtJ0yImF1cnHGeK28
G5+o8kayBluS83yQFAt2T3nm0uMGAx+Ps6Z0PWGbaDZBEqeRWJcaeoczRD7S3SQk4a0Jq7OPfptP
BvNK7ZLCY8oBpcibqfNe1bHMsy/0oLCcy8vz+aprc76NaamQMehQ7fzHAZ7LhT4pZj262wI7r/GU
/kBWO5dpUKGGQdIwvcrkogyuYl25W9cwS18ZHSeqcnS1lLtmqueBOuHIc9TMA113WW/LA7cfBRgy
ainOI7k5LFf77/AkBB82V8D9Cqus3g8yeJgHz7t9wvPVwTBdQgfpLOQ3j8A0uPc+sVDGVnr9FsCb
vZpApuwKEuCXmawbe3bANlswR1iyUYVPHO0oTT6AXk3F/v3h9l6aPaXZKxJZpM5SUSN/wN1xmNM/
G22QrPQQDZ9xiitBrAoMbmoT+s6MuoXltObHlR6uQek4g2VsDnU+W04uxJzSk1b3GSoJQJqgN6YN
SziCqHNRjAPHZiqMIDLzr/H/2Wkb7S8vXqzXBiYAepU4+9/oH2kb1YsiOv7DvTEzyDPjYSNt7ehH
H9j1Eckv7QmOqU20n0YImyh/tVAQ68gX/sLrjB3jc/nzEWhxB2Agh8WErTCGM3gMQ04iUBpt4jdn
mXdisn8OjGrfq1UVp6abXSgYyRpAAseHpAjvwxUbYeapmc4Yp0p21aX+e3k3NmVaJfQWydYRYsyp
P53l8JXZZ4kBBT35riknnIrji36dXRaVl5m4UkDtja0zobrQDixa3M5SmCh6Ant+SEaTeQPKkTrk
kZEkUYDPEWxnnj/w4pNhgsOvsjqpaKArvq0jCXlJlAXvN9QYpk1HyITgYpmNALk2OoCHozWr0U9p
Qn4J4LMhls3IDbxKR7OTL7qKgexbzOhs6oS860AOwn13CTZwSLZqbcuce/Dk/xWtmKYEzbvbao2V
UmZjhlzrKLVs4+05k3zUQxmHylYbmkjXsTlLhXeMb1bg5FreU8cfRxVWyCID0W7eKd6Ic81t/+JA
+ENDLRMYYs09iH5SMw4G+NFQ6K23xO773Ucu6Log12TtGXpIWLXbTZGHZzMAyaPB09ppPMs60Lb8
QXX7NMXZfUkeJBzz1qZgOFFjChwIklHaCtgBLSKQaXBQYdhE8+MgMIH3FEIn8l4zddyWbShGyA40
jVWBTE7/nnYcEQ9W7Iz4qaT/PDCwWsZx+cYLDoyTcWn1+JsllRKCZNGOEHQPC90k7X0reouRxAUD
uMjEqeWuVoMtfGyWdEMpyWV8KdtM7Z94VxUPMNTLgrvagOOi+3W9flTk2/zyLh2s/OS2HKpPgMpv
62/uVTAStGyKC+vX4wSluAZqot/c+VmbfvBX8+6NH5twl45DleTjjE7ggrtmzefVueQnIZy02d3T
Pve1scYuRVS3OHBjHlfmwla0bWoesIdcYJs/0K2tlxQIijVTv/Oz6fxREr9Hu+OExqls/Yl9NkUZ
FI9JNbxUbYLatwSIa+T+IuU63A2IgY9uwpm6JW/rYXAiy83emZvw6Idbdk0g+UdwOJvE2BS9isIu
XoHrxg87RhJf8iBgrwWUN/7Ls6aGWKmxfDvI/dnPAKhI/n3QwOmbTb2YYhw1SpAqmQVpBHxYqDK4
Td8pEZBEZtYTryFemEZrhdB7vFY7X5KFCAiG2GWmBm4+3rWwQziei5FGaHV/nKY4y2MDB93pcJa0
Eyo5M3SvP/g8Kp0+Nb3ZdkJ+1927mW7ZmXKsD3uPxjxg4/XSTRQj9B9sHNZuytrS0JBfAAv13zkK
myan5eZKEIA3ib+TFrsMtq+HnM2aOO+RJjgkL4laTftXkjmogsqPdk3KcUKJIj79/7KIeVNJLcha
S2yu9ceRQxsSzfE3GXYjg9UDE4Wa8xbpHsw3DlHGH8nrJ7b15neFk+5PGQb+wCTh/OJMl6kjH0Uw
Yjc5lVdEa1tZKEk5rZeZH2eYhBoOgw1pW+zgfxhO5L5QGU2veSyTP017tbupIT5hoAi8QtxH5Zsd
/ea9a0hQ/wQgKDlGJlUYHKTB6nX3Wup9Kxgb3c9Esb92zhIVZMI66VEeqqCKba+T5OnX9UxZ/h2Q
h8+1FD15venS217ZP3oto/1PowyCf6XQ/QrzH1co5JVruwDMOVzuj3mkxbBz+gurxFcGyHVgS0Dk
v6n+e5EprsMnzzjh3VTxVZbp6IXo0+AXZkDZKJ36h6CGZfmD6OVaV23AqwaZdga4r9Hn8d3mgd4L
ilscUBR+9Oc4EfrfZ2uM3NxwU18Kp9BvEAXkfpmdnhHIgUbqhLQUlo0mfE8eFxDVKlYotjK9hXUs
L/5funf6Jzn3YfepVFcTO9oUuvPWNf7rNmYRG4nFiUFcDpJu8REJUiiosgz0EyAUYp/XariZYui6
Ayqab7Z8ogzgnhD0AmTERXjMKwbjnS90H81VcSraEphwJouinGvzlqLnDr+E1aOGwF+r7vTli0DL
jEv2QivBP82RjCGPPumVOy1yxX5WjN2uFD/LUKWMmdfihCZ4u3OEmqRLSmiZmRg0H8YA2ccmmjYr
sYum4j8H3VZV94mbzCmP1G8YWDA5PQc+MKo9JVLDM8j0ApXY3Zv8OBgAOw8AU0hJkYC1d7S+cd2d
T4TbuJ65rEg35qQ79gZDvRpURQof2z2SLrZkABWNNuvdiONzbT5p7bv4VsaCppfqDCikb2i0Rgtf
x6uV8vVuUfdGCZbz5qBP2Sw7+OWLZEoLpRo56buEw2zGcFKK3xgELhRUZfrH4QbWH+5mPv5Qy8aG
cEFDAz4QPpc+qtn467BEWPJRgQ2ASgi8VcPrEG55FCYYoc2KIN92NIdXQqK0DWTwB0WaH+2lt2C2
Z3YQfezjhVvpQ/ZvyIIh7PWbcaFUpRJkJW6vwPURJpmH6cwdiSg3jxTehgZ14uY6EXQU3rZ/w8Xi
3yX/BAYdqYk6JTbLW9cWACsEEpKnEW7cfvYwr+3RZiXy3P02RBI2P5+ZEAHurMOfynaj30Rv6q6w
Q/GvqVNAyoKo0WxuzIO3A0RTZYKOqzc5On29q0nwGcBKkLi7zGtViAl9x3XMy1OZOI+W2xeXMeBS
hXP0TMguLV8/Ac097JSlXKSCPlmOdy3YcDFhNdhQQ2K41+N9SSRCwKNKNoybQ2nGmCHA0fuy6Qav
lfVhYNKwwCTMBj+xbHisr0G8Z2Ay50jaKEXo2hKlINvVIKk9oB71OjphrhnUORyA2afRGJr1T+SL
1T8NhrR7PIN3K+hbWSaSj54HRqe8T5456Qhn6lPDjFunQU9F8jInuRKkxfGK1VFp3HGd/M6OB1EP
fEV5rRNXpBiw8EUrklsRGWO3uMAmUZkcpBxGGLztTg8LkRkNceFmpx49LEuyByO2/h82M0iRv678
Ykujt7AU2o7Gy+BNFFmpzeQ0b/3lpiG5ZkiH0rsuTPshcCDwYujtLiSg4i4XiobzyMT5o1KB98FU
BGoDiyXPKAykqyzgSAU0sd5cPeguXDAE+wUKdSfCds4RoXn1V3FNQ2nIgLmzMY5UWeFS0fKySsv0
MfwRGSsZ+UZTMxhf7DZDYAPI3Ez8LaIOYWP4HwYXjjNEVDLZBjn8eMjo5oPJH/DJo7AUgvJtmiDa
DkUDNGZfa3kX8PCUOUNttrQl660E4JHJk6RCvyw/N3niV6W8beDSey193fkwnL947QtNHGx5yAIV
R+RqGu5WI0+lzNliZQNCObpgmEkPgMMiDA3L0LQalGdwMRs2lzwVw+401Ov1yRck7r3pjJlnKsY4
U3XU2AeC6uTZ6KLsOSbF37we99D26o/L5chme1VuUrXe4cVN0LyjA4Vl+q5DYB+DxBI7TlXuudYd
AQwuLM55BZnGKCPzEueEW3Nk83XdWofuXhDuGgGC2mgGwkwk7dtxQ3hf8SFQrtK1AmvOv0Q06YTb
hUUuwnninyyKkOiof/Gmccoqgqrgd/5RYJzUEGLepyBNd/lLjyZEFG3vlqoDe6WeTc1Nn3Jj6nuo
IotthXjCi2d8xb7irxWGM7tKvnV7MdYJUqi4FYLbbSoMmmttUj/VIxZe64PeqtYUloSn7RuCU72x
iU10AKispTPAD5wFHOBFQXkm1UlZPl1CssHotD8YFi+tv5WAgiYtckcjfR72wkhrcnLJEM+AWIGz
Z1qrynqu39w9zd2pefKSJhxXgnIVc9oRL0HujaScJRZIglKLvu1KapwHQ/62quiVZqWCGI+K5K7+
1sQn9wyf4A59r5gfj1W1heVsoPv2qxK+HHHJlOmcnw4bGJViFB11kN/cerq3g4QIjynFIt9yHz8R
Qw2RqASRmGxABstBTwc3+HV6sbif3sNjMpvzdqFZbi36QJK8i2kXFe6+/Y+avxOvk+8zoM3sXnpf
/z1spDe9DMtV0mQIU68+XOLSEDo1ecV1hFfx0yie3ieyX8I1xPtLPem0zKGJdL1eqhuy/qG3g2Ou
6KqSMzXw7kTd7wpWbd0hm0+6akmF/LsckYIw26ndtsIG3eV6hltJGFmNKf1jx/6q+59Jv2FNZ2sJ
nrWJpi3Z1oYskfFRBNktb86toYqbhrVzasVB28ou2STsKMkwO8w4BzO2X2Tp1HUGP6bjX/Qk9xQN
Izob3ioPhYDr9fJg7hhy9I5bygz5t+PW0NfsH+XSFpTVLO1m7cj8O6HUfyJLYeMGdITeHLfyPYz6
KW+1jlRGqiStCuDAO2bXRPApG1Liv2SLjs1C3xhoT7aSN7EXo+oVTY2GTupdoRNvtrodr/1tHNSc
kvR08fdJr6q13XUfYd7y9Asu+OiaUNFZSA1HtbBH2AIbvuogB/B3xZ+XGGrjrPwCnBWq9o0WzhhH
KpmNgVWLF5MxDsWEAhVt4H8tNeW0PdIf6AZquFkYl6OrgtP/a1aMxp2asZRYD2KuxXmt3miS5z1E
cy3E/Z9v8ZCirkOC8lsE9XfRfgYKEKU/qf+rIgb4iG4/QW8f4PQeDYmFajfAF3v6CApZmc036ghU
F6sh5A1BfJXe16M2M/w+Jo8qjyEmmsI8Q8heHQ91ZAgYCUXzKtWsZJhFp68c5wV03+rZD/7ub4bg
wu25bmXpTRgTN6DXMYx1mRLr+fpSYGFlZKRvfEMorAyhmn+O2OOe/BensR+mzQSku9d0Aga8J+Fl
SoTawFgqu7z7m9NKw2W9y+Mbpa+AD6RjwZHsq+5Z5YSQa4RrL7PlphS5ecJ40ovxCW9G6Q31fNmS
EWCzwRVg04UPqBQTMfQB+qDvUD6a2JT95n8ds7Iu02WToOBGZMEiwq+hyufNW5A8TEo40bd8MiVe
WxbbdwasgoiqnlDBIvSILGWVvU+51OEb3vP1P4GC6GwqVGUnmbCdRpPdoj+UzT2rY8JmEQ5P1YEY
nPPH0MvggVuUgJqvCKJrs9iYTjnW6QAvQrd3pHPbQH419rVsFgC/FFaK2V7Tip/qU29ZN2Phr8/V
tNVx+ECNNypTs3KTAzhGG66KW2tmBIa8SVdosbsOVnIv43+NY508+33t8ZDfe9OZhzHaSsAA1GO0
RAl8LwBAApZmUs1/+p4RoXpIs/WTMQwUUl2c9lzkAjXsUq61I4uIUzDVRSgZ4GGth/Dp7SRMWncz
Wtufk0ygsOIzK0IeJDXMAn0bCUSVJvLYA549gLY0t+Qxs58Fmlq3NTepDOt2dbH5yju2Q63b5uJM
ibnju0KYmI+lxUpuWhufZyEwLphsw9ZewFL4dyqtQ0alrwFsK8Ch9Lk+pc43qmQc9F78dVKVZxr7
zfJ7RSy9zYGZUrP7gRnDrY43LsCNB5jfM+w2NPmfyNejN92tSUl0OJ8VEfDTS/ROi6cV2c9CjxSm
xzwSQnkr5PEe7P663El/G/07gHzw0F4wwcW5CtlJrzMwGAjw7H/IWTNs0FQpr8C1uhWe/u/T3Nlq
WUr/Yuf50ZTy8z7pMqzVInevAycWRn2p5CfzmLy4rXvZ4yOgEn8WGorm1KwcO5hf/qY2J83PzMIw
S9rFdgJKmvdfCs8lL/xa7TwBWwhh0d8uWZ4/IsuVb0mk99uAqNy5EADXcPwnOQbdWrWU5fwvme3/
e1zkn8ly+OJGLNmU+ZcZMFvjhk9eIMPtBKeLDjpwZGfesVJfJaKy4Uk9llU94UlN+3C+KnZ7D3Kn
QXzr8IV5Km5nY3c6/qNiz2k69zW656lC7CPK7SPd9r6frc/oAP0CgpAYAFAMhMOB2oKKbdmrHpde
0ZidXVLsbTFnn8pbwCTrKPXcHGADDwHDmquW+qZT0qtPl1Xpy46ZqrNyvl4Ilmhe4P3xd9BiP/7k
b1gHv2lvUTmDGKD/F6E3tSR1UHuRWwLh1fGmkBzwOLu8Omzvm2XFSdHod1v0T0HsT/NlKm9mDyL3
xCl2lRssdpGc4ODSlMdhohnK582tTMJaJTQ+zXlpj7u8rvseneUjt/ElTUW9bwAhdPXYc2/mUJLd
oozwJWLrC6Hb8WpJiLemAlUtTv/wa/W2pTHns06hLJzZAz48DO/nl1YWx9ku7sF8ZP9U5s8vOxVt
jpsUxM+FGG2YBFNUUgz0tUQllP7+Jp+wo6aiOrYtTc21Lo2m6ePhEuJ/zoGmcI40wu7NFcm/2gy+
nMu9uz0b7AN+/AVX0wg8UELDiCCzJJnCzZ9TjiYHuQWrod0uibU8I1mM1Ad32p90f1eSQNc04GiX
lDk/zBMpO/k6RF9vvsAz8SRwzd+bD1kHmkVkoJhFCnrQlC+9xoHwfpIU3/yxYMtCKh1VGV5osnm8
KYoyTWVjqcrKtDTzGfWzBQmpyCTkxJNr/5yTE5MPuur/Ggl9w7AZq9W/9O1NHh5oLPnAbcHD2XHG
y7yE8+hM2Hvo106QRV6HpiZhCc8kGAq3xhP3pTyft8RzF6yAvxbK0gB1yTVxJaeL81kkzXoqC23+
FjKY9JIPJrfH5vcJ7iuohHo+cB4oj+ArisH67brqZAf0eviV01m1o4vlr2c93LAtJW7iBSIHeV7x
ifvMBFGnEStCRtI6kwwNGJsUBwjhEDcVj/FkYVtPsbppFM9aWx4KSZCLKCu5ZqM3vEifFHkifil0
rwM3Rk6n/zdbQ1KK0VhV6zLXgXqa4voGQonu/+9zutZX7Xc4UuU18RUsbAdiFasryQ01+9msf0rp
UKmYfyvEvqW4tEXjj9NHRgGsPqMS/3+BUemEzt1vlx1oR4NGfiv8PGmKDjPqNSGFsi+s7I8hZ7Ae
j5YJ7AprLHBFUYc0octCyThj0RJwAcQWwTeCCa84By20BgY0iLBPEWgP23OgX1NrF7qJWZNEs3MS
+3ospG4nTcuVYxEnXJe0/7rROm8SG7kMd5hdcAhka2RoeUu9oA9/Jmtv9ys7HDn/gNY8gt/1gUgp
pf3x498zAoib568P7hGY5b9y2gyQJZOI5NBFRHqLRC7iPtXq4iw4ZL1co1NMGhK2pU54uSgpy17Z
oI7kT8caKhDh3w617Ftogy5ZmCcDdVYeLb4s+3ZGVcDWfFAINmyVbnkinbfSAXt0P9iJ0QD6z91W
a+6oj5OSiyPUuk8Xm/2vSMx1iZYEkUmWwzMZoF8L+bBvJIykDuQXDRsSedh1WO3hvIiUtB0eNOju
c4Xh5mYmAQk1fw/PB2YQz5BKmcverkh8wB3D7CIrR5fdOf20UHl+cLqrUUyb7chX+4F/5W2GL48A
lithi6SazzYgrCEidzlwowlHdzcB36+B7WfhyrHx42pUpDTEMx78m0oVrPcHrO2qV5dtupzbMfnC
mHI4G1fD8TrGuAGkNYUADDCNkQgytImWEsxYPqrRelfHUQ8ZX10b86tQ/0XPfzcnWEMoEIQyPbKn
WvPONGraSbTpntnP7JOhjJ/6auaR1X7afzKb+sm9vKuirDneO7PSrw1LPCEmPaT5wCi+74JF2e7i
We4pYWYm45wynWEgduGPJbpCC9A52rhciTTBlwwbc2Dl5PeogiE+82Gk4N0l2R1qVaz01C8JUBHI
BB9CEPovYRDGtgckFB1fM5k83nUJ64Nk2lbTutaGMZZYy2lATRQ8ebQPzG7SLyyKjXVA7FGDTHhx
e+Om/5bjWh068U+Ef+5hgPcfETABTRh7Aq3Qf0GfXRNK+QvOAVGFBSCaV1egJ+R4iPesB4RzHaH3
RdQ12osRTgwK0Tx04sVi17JSq3exqhj77NJToSdct4QxMfuVLRa0xa/XjK4U1lz3M8CQelzY+be1
neDTrCp/NqwOXBk7g8ynfwgjIlZ07kARwOS5FUbz6NngIiWOTXRNI4cyBl5GSMaJAhWGfRkIwhgb
UuSjmIcNcgZDjujYL3svXUxUXycYgseAzXFjpNhQP5RU1byZEzWJwWCjyeuTaE4ebN3aEbBLTOgf
ELpvwZnbVJzzZ89fFP6JYRILl6iBjahoOTwEOw6kx8zRqDJJcSW9UsPuODnfqiHU5WmwQzJ2wGXn
Hr1NgfIflvoCFdxUVYAe5aBiMpo+els8sF72el7JaOyF7jWzU0ftzRylY8WNVWv2gJs35vFSwLv2
Qv5i9LzaX7oHKW1NL7N12zQejT/my1OFodo99J0J7AfSPtA3Oj+tcjEFS/OiXKbnoNg1EZjMnMr8
i+myMW0Aq9oHzCN/ghCQlaY1IQuoSfi0MH3IVpdBLbvWPH98jAMCVSE6surDAoa99cFZvS2LL0b2
KLehEMR9gAcC5NCgfVPAliGbkF4T6BNnsZQt9GmphfIhFY/iovnJ4SQNsGY7zwhgzO1LLu2WJw6R
M9RxWzlH4/0WdfmITtiTCdHkeqNBNm1UdQIQjOXbMZpDSQ6svKWFEmPqtCp+0/yXrshLhIL175GO
UYqMOKYt2LdUQXazP5CF//tjcP+/T/nHxlwSQviXbcP+RWC7fBVwhk/rctPpQtZg/Zp4Sw45jJPA
LrHjub1Tz5WbPZVc6LhN5S7EoGGtoHb1T7gdFNU3PbpY+w0eFhB0045sne0s2+idkokrEOz8ZPMY
o2TiRw8UKfIMq/jZGFwwmfn0VrvUBOXepCbX6miamUum3mt15y2uu4FqQZ/RaSticBbRvMXKVG9t
djQp/bzAgc3sUil2+emzPKZl8fWIOWq2PvPsSrMQZOMRi4UdmzC8dukI/gKoZPR8PGG8+P3AIdct
8xvcHpf+N8dVsTqH4uBi45PFr1QGdzpy0sgRN0fhd7aPV7xOeAczMX30bEsves0qgFsgRXIoadyW
/NeqDoMoh97T6Pn6PCMV4bkcbMHJrfG5O/MRZwY27sQth0kO5ozVmhb5KarWEMHRhUfClLOvYZ/H
T/hjq2gTR7nQEZvcR1oXByVNvuLW3mQ+FbuLs7ismQYm7WsKQtZya+O9VY4X0jIaxVh3Tt8PMzA7
5znJ32Apda6qJH5TV2JBQKeCbvqC/yePK4nihhoLbCJ2H73HburT/ncUWHyX7IJV8F+xWd2z1iyg
3i7nojxIz04TLL8tuETFFBzyi4mfCcEy76kNy1PmBUSwFkq9u2+mSCFEkJPhQMk6CSs1mYX8UlzH
pU6jithD6hRNrm49icjeyxl0ERmIUupOc72fpX4iw56rjJD/uMI0qMgY5e8+ceKF3Nm9uXiPglFz
IjRRfIwzvagORX2KIdTPO3EdogMOz1xuBwLUXuHPikqPMTATL/0IsMH2RwrQVASsk+kuv8wmel8p
dEe0t9j0bYuijceR+B6v32YAL2jRvAUfTCWLMlzVZ3SbYrQd3Xxzxn1ML81sGQgiuKYuywxW7c+M
Azl/vwUTA4Z+l3Gk8zmLXWC7W3yDqgGMjatEiznErOtft/tqMX0gRZFmq8R4T33Yn/ewY1oacvdW
GYqYFcXow6rf+qxJGByvOmI9WRRJtTimVq/rVy+kKZ39ZzJHHavyx9VWHa2dbQfX7DuS4sU9/vkB
9zQN04ShlaYOyOt44XvTs3mXKxbUzt001k5yhk19moXeQLL1S1fxAIQWS+fyd0b3Ea64Hq5dpkIV
e9dGRIQuO//ywBF1xwzp6J+M7rkjiVaLTyIYr5W3GRsKmv9ajZyj/GaqAzM0rAMgUUZVSh+NvGEU
m4aLkzizqNha7DfztQo1IkTyKK2axklRX/1/XKAGpDiy7T7b06JmYyhy2iAiyo9s2fz5XOtnEnCU
TAuuVNagCw6KQZe/EtbsGgHwn5fPUPEoHAC1y7jCX7peLx5wrMb+srMk56Bp9sZdwoDxZV7yvYxG
hzGkA7Fddkf4mRYDuLlz4LstJR79xnevrzug5eqwJBV9XOkwP0tC6MsbPsCKv0TUbK32l34352tM
wQ8I8kQHBF+2fpAkVtPWeHv5VBgi+7fJPU5Tczj0bEYgwRW/XfmEFc7+CQFNIrg1vqBWmwdiaNnL
/550/UdcJvxRj1cxmeKKtc0BC8nipb3bjWDyGQ/hH/t5+3rgSuj5LtTZMfv+uj9p4olJXr2YfY8k
i0rtdlz0mg35y4r7EVILRu0NQ+K1EZpodKW8sywRBl8J+sO0NZobVq9Smn1E7LUhApMr1nGJqQXJ
lWGduAchSwr/+Nh4dxbSUfD18j1lsEKVE+UY0wqpTURMHJNOrePujQG9aCnfgM8DrB4MhdcZGXWw
q+sK4J0x/mJfylIihbHSyMMVUKw00a9TOXmnNayPKNLA9qLbBOkeXbV2LLsMGN1xYvsa2Q2oCblX
ixiD646Jh5IKq8bHPn4voadJZYjKEpR9/scC7L7qEFrUS4mrAJDyO46WRDmxp0VzMxw6/srOuxHG
w1spqGIlefKQgIduLH5XcVO8LCes0CSOPsOXlB0nLnW9EHODfPjS85IB6EGbce62bKHjutiachBf
B4KfquBK2f1uqcaB2bvpVafALWhG5qz1Pm4HyAOwtfQLTe9XSXcVQBuWuJoE5flZi1JzV0urz9Wt
8CDV46+9cMyyXZWtBoYrnFn5QwlVScZNUq3lbKmpfmjrMNr6QQmAKt0vtpesTdfHj9Iod87nGO2v
tguyHY2okxOJ7fdKzbTVgz1w7O6T6wsdb6ABz42VqmmBoN01Rgrdd3RfFdTg1nqeXBJq5q+VspyC
5lcOkMpCrFhCn4bM1EnCFtcVkgZ/FmBsro3HawLiMQ9uty4b6MMnfZ1/1abyFrdAg1MYHjWQwU3g
IBblD5tlwe65j3xJOpC2uSrEwyb91o16j5ibb2XCucELXyOvZEXGVc09wTs/Qtu7bbh1tNB9FRmn
KLQaoMSv0BHktubPMIrbRCoMPwv/KaI+w4xSJZrmPdJZ8t3XkLIAoKvynmZnpD0sZSPnRGzLJ1mg
516UrBjRmp/1XS5XHc4PoUZNXP6Kx6jzRgbWDWxWbilpNSAj9uU+sFRkcDhWcx95Uui5sMcABmE1
vzZSZYU3XY+THiS5jEF/drN7sxgdtwf4TnFk7c8wHATEkAI2PewShght1uPeetVPLn1RQM5LVOKA
ZyD0lc34a/3W0PrvlmeshIYgj8cnOJwNdISQWpFFuKOzGKDremzAangbtl4qGThOIkvFXilHA7y+
pgsTg2+XhL62ZZpqAnusetAEB3drmdx3e+p2jw9iID7Q8CsSI2Ng4tpQaTuZjxnSV5jwnOdejPez
ukOyqC1VUp6FmBZlVBF8mydk1LCOX1RXD3H5NCehCSmXBWoxjTuAQ2eSQrdB2FPa//MZHCZZhZ8r
sMEFwwhsaQEdcu42olXNN//OYcngVOM6IavieFLKDQeI5neQgERNOUBKgPiqeyyuOyerXrkh8qaF
vyK+aSh7PJeUS20k+X+Oq2XIhUM4b7Ttpji8z5Nm+9XECmCyqbaac4Ryq9xI+5kMRllsQfAZrIr/
QE1oL+rXj9m5mwieNQ/5ce3S5EC3jmKwaze++ebhfab8lDC/oiET1a7vGG+U7Wd7U4VbzP4TAEdN
8njyy1T9kRZOcyEtWatpo3iaCnZOwV3E1Jq5BAl+hiy7adXcH3mSVV6cKGOTd/ylPvelQ9YyKhSP
4lsi+gfmkD1leJ8XD/dzagXzZKZLEwj2GNpV5HzalReE7dwsPcPUpMdbFVWWHdjYXRqBVbjRD1QR
gA57P0Vz9CPJGgskSzNPthF+u/wxm7DVYREwFa5ytCi2TGF7KrDBq4G+S574NY8PvsK3CylY62MS
QLKe8ffATp8dNp3MtlPREZAykEOojvN1AqLpeGdJElpXdHJNwUzOY66iOrzIX3X76oYjkugUF8hO
ajeISY8c8UgX0go/KgApwC1lJKcFihzMSsWwVhWMIx3tNS3KWiomqS+SAZs9YaoQf3WSEpk8nVF3
jJag8cLebyJrk4CEX0O1E7JR3o6daDjCBU+VTGMvpqb/SEe5ayIS3YAN3LkJQiyOdAuKqjO6qVGj
pDvRRVye0jw05z2nBdvrilzqpZN0AJ1ETxkr1B8+gnTYjopY0CJxR4EoP+tF3FshpDE5/Ktf2BxU
opeWhlARF2/H9FceWS/c6zE7GqcUtLtS5Vf6tvRxZShZVwiSX9xr8k/McOi8hp2h9xNaKeqHV5ej
7H1Nb+top8pf9y8esM2Woy/lTO8DJgBQqVQ5vYrlNNT+8YivC89fd12KkBpev4h//Xs3f5DCC5K0
D/lmLQLlvGnCHOvd5kFKwqDXvixzyMUj/4EUr1KaWooNFsu2JUntpFUXK5HSojIZbcZAejoMK8oj
1byIJdn3jgRedqEvU6TD2exYgDIp+YOnK8UuQpzb5dvjQuejkkMJhziavA4/vLOCz7ms2FBmuSM5
rVYxqU+WQhlffn65OAxuPjcfnxzgy7vp4eKjJI/fxQOS8TjGz6SEe47O2RFv/e3j6ZpcEu6kdfe2
6ynu2ghbFE7CuqRffcC1MItDitOQbcwRDx2iBosXz+6KiJnNjXA/5isdpCnvvOQLMEnP3MWPh1v3
d3PB0srP7yf6xk7q7MSyPL1RC/6NaUBJ9BJDsLw5GXM0rPiXehMdSFkkc5Uk369/sCzsMpsLz2pJ
RTKxwplsuA5ljJLHnWkDF9gIhJr7aYCQAz2wVCD9SlBkt/U5FpCKTHypzgZUBqVoaTscQqUmWvUY
7N3+As/cd7ijRewaNoRQEcT7tYtMHi5B9zv4RF6ZTeh0yhHZ3UEMF6EIh8w1AAFEsBv3L52oyYP4
dp9wUFn04n8J2A1j1fZkLcCg3qOhCnEru6VodxtY0P9Z6yl8JnEXJkSzZNXXo2RF3Z4vJ7fCzLFh
ANzJIRFr7+dykkOXh9Tn9iaqoiksbKBuriSeosJrZDyI3td40ZsqaRwXz/5sSW4nT3N3DVofBsbI
cp0BYxI7OF/eP5hAamcMt5GkVxy9W9i6KwYg5xYWa3GlNsThSJijd1j6brwiy75+6KNMO2BiuYQA
URDXVzAFZii0TN1cGqAzQ2DQ/DgEMcHfmVhogbN+aTvZEwGR4yVWVtD8kMREIEEN4tP4N5U9F4eU
IHDegyn7MGsWm0nvp2cQ0muMWJnJP/ZuwAMb2PAJstG1niwM/MUCPkPYXc/G3rWbpzYRmXaYll/V
u+EE9sv/xD9K0z9dQcdEjwhXgZEvCxDv3s1o4Q8s0iOCKdaIRBiG3Or2UFmDu27zHFHP49dbbvgH
AkwYC8lXpi5XZOcf8+Jo9nHp6QyFWBTaApzCBvR4daRwo5+PjuwNyy7PmF+Ch9MbXid2RTxdHrfO
O7cQENmLRSXXFggId0RMO/F2sD1G+7+OtTv66To2BDrMwc/LWVYy4RVKZJgoFtO4B8kIT4kk/Mep
Z6IGs3zTOyQzrms2T1Rg9vUguUggHY/QiNQhpm8Ft9LD7bpV5AA319XRtVWNPbzd7kZu/gtKjrOE
fmVgO1gw2oIuF/rYoO2lwDUVbbaSyZKXebzYf/Gsm4kxBiXtnMv8PX81rhaTSva7EXGJGw/4Zklp
ldKQcs1nHinC7Da5Oa16knGsvsVBdvJbFXZE5JSgGX755ckBXye0/EkSH17FJ6wq6AdpTWrV2oEy
TDXwQz5IpGypqkPe7E4a3CvPgAjtc227IO3Eq9l+xwPZQWe/s6ZQRqocAt5wtgrp+p9ie447RePW
IWOix5XZG612A5uNjFkXKdNtW8s1fQ8aqc5DTuXLDQqtdThmyom8VfhzLq8/qptFjZCvyGo2mE/Z
jmOH7WdW0yQoob26i8fOw/D4vPX5StVwrZY8lRs+GC43g9wUJ8b/tU4KWPga+srdidlCFVcRjP6/
CW8bsAmxwpvlX6nvOYI8o9E+QtSutg5RwKtfT6YfGXEpQsoPQ/vVFf7PxbdR9J/bpPc5fPSGEjaM
Nx5WuYtdl0AatgpeqOapgHJjtO4gYRDF8KqMmWDDdMPc4WoJEQFsg2aqT6wf8U6AdJb0XMfT1cXx
0qvyeZSM3KwChq+9N5WZ6UuViINN6jNeItsSLFrfesh/vHcWaZ/T+mjmlsR5s2/kBWTwwZ+vrEUr
N76c3lv+QaGkTSj6Yem44Jwbf5W4D5Q2DPp0M7TUUF4EAYNFJH61SiMZeCtSA8lXyj9Ftcy0RE8a
d0IL27gMhM/0MYhIBzVBJoU592YnMrt7NcyB/hpklcevGNRs0Suzw89Cp8y1qLZcuyapuDv3AQc1
Dqur25h+MR9VdeNWq5/2bPP8DuxPTpEHF6pyI5QWHDouCC3ns7NGpaf7h0PbFwVDK6nKDlaWv4ab
4m8E2jB384mBBCre3arHuZSCBWo9PGJ2KoVYFUaZo6LR/adb4amcRh/nAbL8OeiCermofu6pG+hp
0hR6bMaJqqrh9I1oEf3b4svYrM/llM9Neav/snBqUBeVfgTY2J1oukg+9E5ZjvqMJbuutC+WO1pi
7qPmVGi3bTOY+pQotmJaBsOxKJieybjJFlXHOcMJRDeaRi95tFJRqvWB+2kNsn1u7zijH3JRjTA9
KW2wHK0e0I1YTwjFJIdfwq92QyOIz+G9w9hvtujnkgTa+rWAK36RS5M2BTZmeev4tz21radZltk9
QnlX4CmnFcTb3RXmxNVWXodziWLYCvgKMUQz4ggCsdajEMF6IPhMIzX+zhaqkzLeyLAE+Zbst1OX
8QpuIDr7AoIn2h2AK/Mtd11LDdjBsHFKmlQrGDN6Gt3mJQ+WVUZCJPeWXqLCEUkBntrip/Val8kE
ESKR0bLYxjXnn+FwmPOFOwa2F2AgZMOhEirDWfPpyToisx1y6jv7KVqXrzLLOe3o4wFwOhTPvsVY
5rix1nMyA8HYgBxviH9Nobc44TOecSwKIBfwlV6ydP1Jxnge9gMh6DPzN6PxAzymJz/bCiI2MqHt
J45oWxQj2P1i/2IDFNAnwE9mnrhA9QoEy7oMYrVcBkl5991IN/TX3DwB0BwX6vcPm6XoV4/KeZiL
jISCtjJOKGyANHbX4cbaCFZTiAOJtpd3qXHoYbxHn83zzcy2XvT4fcAPUFrFLZ1z1/lZJcCm0vYl
iqPLF7Ke3rizQ38g89RJok6/aS9+aclNoSJuWXuxZWLKGEsaaavGCRxfEYjAb3RydTjlfO20ulQF
3cGsLp4uqpQV381NhZ9+A7YFXAgu6HxMduo3nR1nQTkJ3JtEogO6lylMe1rRZxTnkcziQOU0B38f
x1hCMW8dc8O/WRMFO+Uy3y0TVC2di4c1h/GCNWGer15GU4X/a7W31jzETe0JkKxRUzyPZqHntWB2
hYCfCtydgOc41BQu+8thZLKC7p/LdZvUus0eWJU+OTj7MvEc0r2dN4R4Gp4Ud68NRVLR0QLgr6f3
fyYDSRoUrgKK2bpQ2rYMoUC8UrmyuvnJfMggpSSMrz/qM73VMZ3fdR1GuIWtcg7AWm9rbcf0OqcB
pNK/hMvD5Cu+6VmDhKILzICXUtse+7yNh8uqa+lp45qwxub28c1OtvCDCtWtfma3l9wlL8y4ZpPy
kxXFkp0kFfr1bWteEum0gnP92vDJAUop4wqxQNsEivKW60FEHFwRqTUlFxM2EZ9eYCraEBaz443W
EExyZRXiQS+3GOflJDnPf//lRz91KyyitqPLQqc9PQMhtOA/ogaO7cm/MajitSPl9h381y/P7OlH
23w+mxnwwoDb7WpiAh2HHFjU+XH34JDSBpQm5iJx4qtTaEYI3WsQlJbp1z7dZkiQeTOnRpSqRtWV
n6uap0j5q5au3NuUqhpgw/ySMZIo8LfcXGGs5pw8x9PNkNXdWi9Rcy1s1A3HdndrvEcRGdVgicDU
gzMRJGBTZ2RS999R6/iNgpOC4T5dBDDk86J8Ql4TylJ52lVKC3QgN2zEQje9tFz19hlITvIQuaGm
/HgnKvMyp+RgaKV0yAXcL47hC1+FFQOeTzndibZiN2Kjct5WhYaspDSjNih2GRqwmY+9WLgU6fWS
Idxpk+C6RGSimOEjjH3V+rj2Si7v2MOKqmonBnnCEnyBIUtikLtuRMxSR+ni6VK+KDougjcteZAr
QA0b9MxDmSz+t7c2VEraFU9nALwNInOcAr/vPbyc8aU99Ghk1IWc9BKdIAdOyN1imy4ZVQ/jibS7
q49KwgfsSA8XXYd62hjANVtn5libR6KDDHRdKYEPdPf8XRXDAJ26yeFbv0d1tuMabK2Vm2swY+x+
ciFQOxjoAcpBgsHq1n/gqkbv6vvTX0cj7+oGPwctGN/Yh3qwx4yWeLXYD4Aa2Z6TYkbp4xnJcRQe
gZWzRmp0mVxYHItUY7HY3feAvJ4IhAJ1iUtlVisw/Lc95z12lF7V5l1fQR/ifZMgaEfu0ecJ25eg
2t0Cgr6F+svzyzfuwQMhvC4fayEJhjVQ9RI4tQetu8WEzIGsG1IeylgixD7pNXotWB7MLnmgwx/1
f2pgwhqNt/ew396cIccMW8PsXhy6t0GvqVi35RoUq9N8n6vtLLmQJ+NU4fvDsxb3WFUqJ0QqnPe2
a7xyg4ASdK/H8YnFuynPG6XEag2bHX3YHuqO86MLGRd9VxUEseQpVSXODiBJS6FcPGlGlsPCX6QD
L4k2v9GlUEunYrZNqyPsNjBBoH7mp8zjpSvtH5NZG0tHDl1rRGsz18ifN7GSWX4dyNELIU9YgBLb
LIvPIEQOpDJ5PuTtfsoR50Yr777Xvc+fEE2PKLxHwhGWMlaoEumsMqwvqP9jF8i69pAjmcsVF7pv
i13vACninTYBFK/sSwbi+IGHthG6UC8eGUN4tIB+KpxpC6HKK+6kGrO8s3s2yDxXWUgqap3rmFFw
LrgLHRKp6tS/HW5bFs6KRpsRgfXIs5Ly7yTW1z9aC62xUH0Y2RPxnmYNaYx5yTbXlrK7+XvK7UZ8
R+Kq/3gHDf+QTZjAr+YloHKBDp78bj2eR0yA7UPGD8Mdcb7uNpm2S747Kz34JEXSu0AGqxkwdASk
2X3Hqp5xylcuIdj2o2cCfhz640zpHcGFemJQD4cFfjvXYmvnXWRFsxkKygeqy8LmMKIoanUqEwzT
xxDa39QRT8XnsFq7i2ZD+GYCLKr5sNWvPCxKIR7VUjJLnZjWtuMqwSTAoQahfBiAG7TfOXrCQ8M6
Am7qtsmMgZtPG071Hkmn7xq/ROGxSsbjXmZ2b7BAD6kkb3ndHgo+FCXLzntZ7R+uzAty3jupmmH0
g3Wd0vzDTchS07ltDI2ymKzv33gG+/7haZhJjlNFGgeUWli/fflEmR/FglRP8omATbvYk9Qdde8t
jmvXZGG2sdvNmy1QP37GzUhS7Ib+B59OQxVDlw9fA86rkchnU2Wh4ZZ6E3RpYsF9qN8yY0zrfZPQ
6bjxpNdu4Ge8G72Bcb+s7kIIseg30T7aPoylBd+UmVjNSpi2D/Rx71U1s4BHz/7hsowevKLeLe02
HFDxFIkuk2si9CA6eHXwep66W3Gb/TBPPmADGILvPNTkNVo0KCP9t9Trr+dFXeUaLB7SAzcX/l9Q
Nd8C7i6myfECXwM/CdQG3JdKvI/2/pGgdnHLHfvJfiNV8EkdJJ+UZJcB4eC8ybUZurCQrkgNNFeC
62Oj7AGHpjaEaTQeeoDRfW4iA7A/eA8qUKF5XuaF8JrhPtAOZio2Vvq80GU8ziHdgQVCan1GGVkm
t0Gvs9DnlMvbvi3QahxE3seEVVSGIJ7+g1iWg1iTcwgxMmbH5/QZ8YtEYbSs0/c6En92H2dOvQHn
IcwXZHwVbbK7qB+JNgzIkknLPun362elTKWVkPfjZOfme5jNaATmioOh+W7KDK0M5/JsYb+sakoe
efuOs1AnPHVJeRSfCkgxoy3QddjVl7ZbasHBp/jVPEtMMXqLJ5nxMLPkm1Gi/nA6k4uCEgVHyEEI
O7jfnryZYPGEC51Ndf3muMS5+x5y2IA5wHz3xbzew+c/xHKC9lk9RsZE5MK/XwN22w6vGtJzqZdN
4fUg/mBoOw8sufhRgQk90iyEfd8df9Nb+9nxcN5GE9m+ZAQ0soB8Q0dubM5Trsw0CZd3lOBIuGtw
zQd0Ha9pjW17jvnvypNBaz+0aZ5IRkT6EcpOWCJLXk11nWCJAAXFd207RhNLutIZTOWZlWeZQReJ
KkPMQpneOeRabgZ1+LgTUxOs/Z4M8otqktdmW3nl0nAfihf84V4ocFpgT2+WEvwTsDifzVW87uQE
RPSrOhs5Rf0MIvohKUQeyJ0Jt8lPLBLcoDx8iWlzI8cQoriEVv1Q067pdMH1DBq/JzUUz3mWHLvv
zDVNhSzuIFmCtrIc8MBqchLJlkgQyjohSh71xPWaAMa/CTc8POO0Pc0ZGWgs7+rGgFrSpY7ngTdT
GSHTv189tfV+EixojeZCMKI6phNYlDcVTyZr0z7gwb72ZPvk1mo3lhfd2L+ryE7m9BZ+P9Xc2n5E
LlFgeapW8Y6icZsUEpSmT/UynWd/UOicu4NgKX9DKeoL4pTO6Kh/jYpLc2lewaDJNswoMhLME065
+28bZwQ7Qj4BSMLaR8raHIg/QuetH5mUqp8txItrvYAxzryeGxTaH6EN1k/5ZSdBkfYfkDhaf4Pe
b4CRaN+MLaN7zVSd/DKmD1nkolwBC6NyUeza+eXmYWe1XKQGmx6C0HsLufyT3N3/ySlukZE1lE9r
M9alArVpdIuYdd/SjZuA9Cw10jJoZOiQmqh3u9qeHOYwmqmOMT7kxUZ7BW4n7yMUuNWWkGZb0xoS
7iELWqmzmju4eHKNSq4ke7B/fxuR59UGK7t7KIi0m3L8xRTQavWdMwfqaUb6Gx4QXgD4wkg/6aNC
vca5FDIQsQfTXJm3ONA2DZtmxWor5b9EtRm1nnKi6a7BYgadYwRqu+hQ4KN9s6DY3iWI+kXk0ZoO
YosOoGm3oZsWfiGBZkGRZX4jlTHtr9w8kr3h+fH+b7CrpeskRJLoVBf/HzKpUDb7Hq4Yjefkxwi4
JGIOw43ZAudeP7WpT6YwsnPywmgTkmKB29Q5gTjFytIR09LW3FCcBdIi5XKGw49AeYlWi40gJ098
P21HRL41zixJKWMMN6jfqOmKc+84zU+xhnF4rcF6T698S/SxQ2uZ4pVZW2oNP+7K5WzimBCdVhNT
X/MqG0slcB89lCIzQrHPn2+wCGamv2Npsr7an94Qph0DAIB69TfxSRK4CjA31zAd5+/xZYDhaF7a
3BOblK+zAfNQ9aJmVWgWSxGjlVR7N3022FujRQMok091RLiRFvbM0LJcYFKgRZPNONAmtr/AE3HX
LAQ1L+T7vfH3PZa5n5Lwkui1Y3aXtDpBD8IxStVSz4kM4lg3smT3zAheNqVm2ZBCtGMTA2U+EB+j
D1DJbLMedxrUeGkrafF3NdkBEV2Cey5D9gePoRbHrQ6tKodizU780lktZwvef4WV2kjqoIyShlu1
jwzd6rCZ7LB1dlDZ50LrKn2gwXw2zVbOzUe5o8MnEAr5t87WXyyVzMX2eeBx9jIN0R3Y2m+hgRj0
M0Npa627bVCyxGfilMBDapvZmvoB34f6C+c9DBGU1DdGw18mXKJxvPmG/s9m7+IrKCioGVoqV+AP
541fVqmFmXJruvFq2ITW+vBhO6n6getocla6bwl0E66d5e8vxVFFMP00OnGt7hlOwKQt99b7M/pN
wWBki5eZ/67ewBWhq/SMPVKgdsZhrwxOU8R6LM+NyUmJTNnxN49plbdsFkUWZkiHh2kOHyTGkTCv
/tCucff2gblGb2h4VPSYeJLOBsjYZwe1JwLki+Kz6nYKAmdBvLtDbXRuQvzuxKTOfIvZJinCoKl5
VzgrtuOCnBc53/a4l00fdJQM4vDiEbd/XIIg0us2vxx3WMEHA7L0XeiDct+dS/LBl7sb8FDiDYCT
aT7O5oWLbXKd1M9+Fb+AhBE9cdIVrkMFmNe//cz80JYNvHmu8gRnfVq89t7f72SA8iYZ35rlAsbD
lDBi/z6pk6WG+Z1IM+RohD/h3EFpoig4CUkNwsWeZlnHxO1jJJRi/p1Gx1IFfHZPxj4RPao9xKwA
q4FFdQoKXkfvXf/FdiNBOUKW4a4hfzzq54+lj9lGTLNjW8kP5/1lI0dDNO2HQaGNpN79Yu2jYj/L
uaFnu0nV1jaYhRi5Pwq3Dq0h5Kklx7AzW7Z/vDvkwpsIV3demg6Gu3jHTkPQktXZcFmrDiz9lbp3
DLtWWwnuEhwddIjhxSi1kYBMcANKzn0zV/GVIovIttCCuUEO6NiRLF1V2798Ao5joK19Kc3/+/tA
px9YXeNp2r892HTt0XCEFVHuXVPoNdkPH0ufOW6juS/FTS4Ahi0B/TRcD4fVk17FynCrTs48Q9xb
BLAiRHwPepo6C2aoNAP2hOUQof+bNfoOW0cvZvmZ+Sg2HhSotiXN4mgmz8ajttAfFQaZfY1ReJ9p
BsHje0MMZGrQpZTDBkrwEfsFOlA7MZB4dMWkG6a/eGPjROuW27SVIJQwzD7XANuGmO5Wh/QLrA2G
ZFIwVT4J6/EEqN73CZOEbam2aK+ftZWLL2gVEnGJ7jn4+e8EozqMSDJ1Rib7+41OBV964DArQwoW
BGLGcS4ZpJAbnokKCJZ46uHYVVg5vYsRMO0lF0UJmvkdGBcVYwe4wgKmNjYmAtdge2PdqRVE97sB
9J4/8IbgoRCVwvMkqv49dKpVx1mq8VqK1MVMdo+P8d6Ymd564EFAQ+VFreij3kt5gX5DavYxFV3m
Py5t0yTfBFDNYjUIW+vFpal/8i/IMDvad5fYQRDJR/JpTiB1nmjvoH/1y0+HsNs7U1YIPuBta+o6
8ES+uj9Sq1Dseu7BpS0q04OQuFH6o1meLAm/wz8BEaB8qZM7VnBNLe8y3OZdMpCQ7AEMsqZ6nhPb
6zRZ/HwCu2B0ssV7Toplll2+m74+K++zQ5c4ELmczCm7XTZfg5AKSz6B/jYelVQM7PJq8p+HWvZE
P8gTQmElL/AxsP6CB6J1exQYanQKX9HN293qgMb5DGnPnwGpY4fcGxj3AR1lKo0apcfXNgcEYwYW
Bn77q6H42kGwy3vmm3CPS7RFNNBHNhrk15TnTT9t89smUc+QDhJf8b/idH9MqQ+tK1t9ZRWkhWxe
Cu6LqfjAXqDcbRYNlu8JB9j+Gui/s0ZY0YxR1g8B5dkr/Hh7mPR1McIoEwHqfnIChUWZjGcjm7Cj
gL47ROSISIwliV9OY8R5iufZzU0sunDWpiSHHXylhAzy9it43LBWOulYE6PSqSdXYMDVqUQjq7EK
dMSA54ousYI+hIcP3roR43JFlg6DOo6aEJclY6luz1kF1yUv7L81+lsaF3fq6/5km4riIOocJNTZ
EadqTzxA8MbfwNsahlHKz646o+4zzNJ8UkUEhvzMcM1qyPU9Y6mUCaMddBlsmUAjrhOqunHZIU7n
aRb5DBh0UQPzzMt4qmQNaLabnQtGCeTGhV4m775DTa0qzc8c6NhJcp64+8OxjwLvxt90yR8y+Xjr
U1iQ3G5E61lVOrS5clnrwyCzlPqqbQHYwWKX763iNa3HvH8+NuteoFdg1bh9JZDhqdGXvP2W6hFF
lXeeh6Mr39Uh0uZonuYE5QCZKLxS3Zojk6yQhGMgRQL5a0YMTqsgOHsxQSQLyua2eG9f+C3u8Ptu
0oA2tygKzbkbvrw0lPeDa289GsP0IayF2PiY35gqlTxetChT7kuusfe4j3RtI92ENhE3toRYkVvC
HxC+7ik9tmtNAcjHbPzqaZnBFVTVzZyRooYiqadj5i1fAg+9oTb7iA55NEPwJ5oJGddWaQAsR3/N
JOBnXaqKWPpB9iVogIABh9M0wxBxpaZzmE9e4vL7Je9Q0d31FuSlGUQjcTacVBQ//9AF8UQJ0lrC
gcbwM0O1FqMVZ02o1kA2xPOJdJCA/rKUBgLiS2rnEf8KjsYfPCsKR2/QDezX0gAYc6rCE0h5TKF4
1QB/Nz9g54YtkVrgqOixjfylG/bx46R/T5oeWGiuplDjPD3AYsphjDEw8lUliaffVocD0AfPTZ0N
CIsF7bCA+8eMffg9TSJLRrqUy2dlM6OSf0TcN9NUUnVT99NAtJaIGrJZWsnOBtyNDVhLal2oHxln
3IxOS3HrZrs8fvoAD7HVbdFpHMXCX+9oRn1tV/YB1U2j+eLtyjO9aTLD372nDYFit8ygN9uUWSZE
x7ymZsqS5V4yBwfQ3R0z4g8enFt54rItmYBrG5tXlj5XnkXA83RP6IodDkUYV/F/95dtI6R6dyig
xiwKHjKx/FSFSNUf5EUBDzSjcPG2z1ZyhVp/e/e0foyldaK3BDNV7kP05TyoSr8s9g6VHjNs9Mx8
eag9/538w5MVqogu/X/RtpgEClqiPl+iI36Hq0T0YIEJCdpyGKlODxiYNwBx+M5XsLGHlRkvlvzL
c4S/M8ZmytcjuwrB6+K4UqnCEl7VCr/XVZ54P8+bHOPu9tEqVDEKHEC/x2R9Jy1uGRBWeG6AqhHL
jTE14y2iALfv2tjbmJ+dohGeqwI7Ss9iGE9v8lKKHRi4Uan4wDM1ArlT/n+SStimERgiQgy2tsFY
Psm64Y7tGYkX8qMYGilDz5ax9kp93fXyJ2ItFT9uiMBFkOMe27cfbEM4XMqF4qQdYtjgc9MNO1Wz
653oNphmQ95hEgxv/8lUNnjHUGZZa45Kuejrp0fbOCEEcIWUoDXSII8ZPSAiVFhnnuv05tthnZbJ
R142zkPdtYaS0TP23c68h7YFSMdCnZ37KE20XZjJXU5wlBXZSHxkVwIl3U4GCjwIyNDvWAw2BXxm
QWE5PqMrObpJmg3+DIlHyGVhFkvacv312DFB0eMFXHP9TXc086t0tzsDbl+jX4WdZfZt/vi5n19c
yLTCyg4CnjIgKW9GlhOOQRuvzinx+4EF7nKaDNEl9viXgdaSxifv7rf5T3NIFBlA6FUOxrZH3AVP
V3ke+7zM2db1kz43oinTnotjSuDME22DnN9Z4qFr59KDZ0LB8ht3RiA3FJfMKIgHtEaV0+pxJdYR
CehLU5O5aDybRUoMBZekHlHGZuWQerLHDQUYj6ADId65j6npLMImg8Per3sxW1vlXj8EKirELjWR
nWKA1ayeQ6uEyriTBMhcdPYaKwxlR3GBmGhKP9lAD+bhTEVc09kjKEyJD5lslyAeGPo7k9GN/TyP
YzRG2U40hhQniF9wt6Bv74e3XRwrKwb1YYj1hJ9eFmGsjRjMsdXCobV1IlzKtjMenXXXSnwpIhxT
jcl46W9fmKopt8k6j2Oxh9lz79GxBGVhe4Y7cgf6f/hJigBn7MFMNvOOKFXTBQQs4wcesrIPLkLM
zsg8BEouj6Ho7Yiq/AyiH9wgxaZgmXDox0AHRB2YGXqHr6mvEzRJ8xZ4By/bhGRH3lz8xPCUu7p1
/ziRdFN8o5vgQFH3Yoj/alPFdcT2xOLWAzDo6hY9zKSLZG4AbMHDNT4Lojg/Iuy/5d2dlvdbn84k
PU+2EohB59vNQtYFlzntIEFFIF5lq7SdXz1s3ij77lK/dxc7wxw3NwCDcUjRzjGdr/U0AqjHx/By
fsj2wHJj1jYm7SN9BjWi89UXoHD83ifN0RLYnX7ttbdiTk5BN6FYjVOo3juc2yL9fyR8AQ4+4R3j
LQGgcNfTjefZu3QAxv2X+WaNExvE/D2Wepy+QpVDhkvq4yX/AeVAPcvYlHN8dQtoFqDdf3g6QPqx
6VqxzK2Rtnt7QiCzePwOHcCs5iC26eV3qdYZE5QJjxLNaCYlDRpmEsDQpUn+pCvOC8lSQMExXuM0
EiMzSh3wDnhm+LdCxDaZx1f+zOQrkg1sKvLCTlaOKUwqDp9OaET/CmBfBeoh3mYpaDA8dLxetKee
Kjor/CacFDVm2cFDt9xPYRMhdQljXOIn839Q4+u+kKdGVV1Z2Z2J9RUtnYk2RpzC2ogJjYOU0Dk6
DfDCNQDP2NLJ31ylhXL3R23j6Jw4T47lZ20Q+W8IU0xbTMp8bDYXJMwj2/8TAhvu2O0WLf8/+PuE
I+qKI5C4dRquns7eSEzfEXOhhyxfDc/IuCqJc6aHBx1ZRHwkVpHOGk9N0ZWHwZ+AULwkJ6FKmZnR
VH+JG5KTdZYReuIo6d5k0cympJTe+SReQh0Fqd5qhimAlURNpcZ9CVw9k4WezX/nxNlDf2bykGwq
EJzkmSuYPATA2AhS/acr4JDgcj4fT9fkwRvpjXKJuKKtmN2KZmh5IpYa8YPhlVubwlE3uF59dLkG
xk8zpMhHpPsf0SrlW7tuLQzJF/24mTZmLDJFmY3wCty1ePbthE21cbrtrNLBE2fTzFrhCSlVNLbW
zMY4ffG0HtmmoV8x5+n63y1ZoZZnTLZnTdmu9QqRKqGJAeu17XTsF4oZX8qH0fI2xjZPyMyrUI/9
6Uhwex7I+ojlc6oRYX5RG91QEkoY5/a76EbcrwrINJ3mcu+cBguwjJHeW6P1jlEl+pdy+5+xwx8Y
E+nMppbgWQ0hKKwe+B3cfR8ZI6TYCO2rfj8HMAzfIJtZS1nxCi9NibU1WHGbZAqzafsWWdKXB8tN
W0b7eumsM0AbELP4EQezPSASSnSZITOGb8f2hj7/fnh647vUq4sJahbiqDj+18Njfb0OqHFrHVPv
zehyW9b2oqB2l5Sv+KvQqYf/MQSZ2/uOo1XxIlAoEfnT1D85aZKDYn4GrFquTZdqLl0QeymmJnth
W6twWQQ+jmIJ49mUnN4nuW6bxkQnk8+/CqbPAR3Dq+78QhRIbX6lP1rmTVrbuEewNRVlT26GNBLj
ZxYQygOadn0qCOSL0uhfR/Y1UGRb4YRBtvwibInltUHDzY37GUlNpKJ1OK+pE8kV6nr+Ogzq8nWS
qCWijngR1pfmA5SAoaf8Lgwlo1B/9qLwVsXLhhviGBFgleSVwOjpoWd91+HoA7xZB6cYPJhlzbbf
v1rKDg4vjezMY9qm200/71SYBCiDPlAi/IpZs2Z3vygINPuYL/gxGQiZU5UKRDv7ZnsjjGAP4YmL
JSZwm8X9IhIFDzYpQFnnT71Z5rGg4Tvpo1DKTk4UBcr1YeumgZFnw9VlavOQQyAlIfA/SeFiaX7c
ifuwkVLcqnY8TteyGZz7MDTFLQqaPfZIdQ5K6GrWiBokcbuwpBKqL/ArcFYvjVDrMXWkUZPIsRhY
C2OvJhgBTik5yDe1+9sdih9VHDj7nvUgiU2Du7iFDkBh0L4Ld0TJVvhzjYojrlp8svsX7wCxCj87
MOKMROfBfgCXFDxFMljeLzWW1tQ1MW96kUfb+FsDbjS08K2YkVEGgky8JZ/29B4X2MvEzwEHX3xS
U0IMAiLeyxSaao+vmbS2c75onPJhn43LxkgN5DNquYdjiz+4CsxNIFppQHMciUD3S6Sr7vaxD8Rz
X14VAemTmC20m5FHwNu8+A1kDvRBd5VgNTbdWhJljoSQ2IU6+QcLh747eEEbVT6PA/f54Zzajy+v
g6ZP+QwbSDJfsiZEgVZpeUO9Ed4IQOKooqzndlc/+g99Nia0KHwdZIWeAO6dK1h+M5icCGlYQVUF
pJKULpxUqnCdHGLOAFM4mYnVhhhbl3qXuRXDLCZ959aWmKfDx0CGlwy/Z/gNbaK/kXAa4zH2xhBh
n5hlkvar8qAIdbtFuzTZxe226uExr6jbjlm8MDY1nGMLCH0gKUnksnak7E2On1mgsCez+Y3x67Bf
Klpj6ooAsufRqNZGH06Uo+XOm8ehibTYhAy4+XLEryYLEnv6UggZOr1CZaYYS/p/DInVn9RTt5CA
L1vbStdUIMzbukxwY+lBr/+ipq/IZpSU+c/dBIvb5FTxnWo1PM589TtG167Dz6ZIiLF8unCqbwFo
2dnOlU5l9fc6PzDbNtQJ32QFuYYZAi/ySrw7Jx7PqU0asr0JjZoeTZ3gSE2A/4MfoT5Iax0bj2XE
Lq8fNT+qQ85V4d4likjSFjQO0pLCwl2ICRieQggcMM9Qpe7WXMzQsm+ujizuiEufdApr7zYIhKBR
a4eO7AkKpfhg5JUY9G94p0Mz9KVG5/G25x2r+W7dP+ef+OwKuFblr8PvRlnZBnmNIwSUQ64+X8bE
RVMH8g8bb2pIjRTDR1juBnspawrIDkWB/aBuB5lxhlMeqRszhHiWosX3rHsc1vNFNQHCrsq4FMZO
GIc+sEYhh1twtM+wpy5dxF5uwNXU75fpXovhWut05cY5wBzTMUWLYl7PdnFbRWtr5wJQknWwg4dG
U6rXfmHPODRRWCgKKJjOKijvxm1SHY1pVqMDXQB642u/m3vLIzEyN+xA3oKKNo1pAt4/vAqFyDxN
tbPQz/gRdqvca8313pVA7xqiQTgVAc+Xp77E6ylqW/3aiTuTAJx93zgyV37M19j1G6aBnaOfa6qY
KirvuMBMRdrbCnV8M7u9BhyqQxcqgJsrYH0jjkBJkSZaCub6617/mY5E5oXU4g06Xnj3Kqj9fbkm
5Zt85HZWbL+XlKF/fh0z7EDhhFLTU4gcKjDnoVRVnaiXV+QQqoXfY9YKMZknhZUnj2BH8WPKzQ45
qltN0mUjVu6FQEd6rtT/cAN3bdoETLOQVnzNvccy/Hjgvj1R91WJ6hTtWZkGFTuxnW1SNuNy5u7g
lNH1ZA0Of6BJZPIiZThGEJIq31kMvVLukMb4EGwLNIPXe1YpEac9OPgj6Z583V/Y8mc0M0mYbkUN
3Mn7rCqn/NX5Ib4nlNHGSxmjuBXAseBaOBxJoMCNokuS1zv0fzxo43zJjBRM6dBUsWPI2qpbB3Nm
Iky6JIJhFeU9310sYo8wp+CK5ngxE5rcubrkEhejnyWYRnE1Kar2REQehQRqnaGzysvgbxHWljht
nU+Cv5z7EUNeMhSh87Mu/zWDVkU8/xSOjh88s/Ke2KfAWRLM4OvdyiuhpkuS8b+4NgXYT4/Jwvjr
qc6zFgGf3ERYzZpklnqFQb2EYjtMaHE9tMVrjrx0C/kI6oOJbDdr7C8nDwpsfrrE5aGXtIQCkyEZ
gI45H74WHpoGTroDPOOIOZ/E7dWTkN+0bGJzB8Wmzs2PvaH+3WZiWYS/cyz45Sbmjhs+Y9ioRyJM
gSGNzDS7OnUzqd9DYJTuqmtvPInGZGeV/xclPuObctTh3JXM+UAvaPLspVrcAH+Phnx51h9S8/tw
j12oACnZvyqPLKZlouZkHoDeq2QIHc5UW7WSYPVKGykW+oIkZ4R5kXEm1vW4rffrj8tniIQ8QPZX
hL9T9sbTsg0110SsYiwUDvOEQ2JCNd+CHpijvhUy4qV3bOoIVzmWIfCR5dQvp1GJP3LEjsEOu63P
A3yWjJJJRc1AzyosTVjEKvLO5g+m9YZFLx3ybkj/Sege5WM+g/FaSi+g++RxaegZznk/lWJ3aKJh
7OpnkNh2Uj2i+QcdCJXj2wBUmSL1mTYjMYRpVMoob/jdKHF6PynQyvYKXGzeRs9tDdoEeSh+FB8e
X32QnvqTfuvRqSBRGBz9P/vOof4wNp2IF7QtqKWIeACUtl0NtBPHrs3XHu3nVjLg0H/ptw2/Jr6U
i0BQhIGXpks2NAg69FAseWLM0+CUxgVRo2QpA2mbm5ThZaPfg336y7Bi+tUyT7SuJeh5ox5s4uB0
7L1VhR3M0j7d6pK/nFwTCXfcohX5f7Zm/hMBT/wTn9DfWKwCiP8z+dzg0hbuoBQua4ifjXn7SCaO
zoSnMFxx55cQXI/btWzgavtzStEjJDh0tqhujP5nvsExNg1rujGZA00UPvGweGO4GXJ+ipMkKbW9
Hx/NzCWVCq7oMsSpyGXzyeaXeZl4OyW7BYo4X5vet0Cxwkse0IhjF+2mpgBzHj4BIvmOnHMlkpHn
RBs1yXA25kcWrTNnGsXiXtmbuz3/Q+KERte7NrSKJMoVBy/21otRBP+ZkclDb6d1Ea1wQf3R6SAZ
CGJxAYBxqslr/WQEs/I1vdqDhtylT9GP7V8E0MiyeQNE32b1jT8miJE39bK3FPY45IJ1BjGMc208
0gw9xmFrVjacXBIrks99X8UrejN1asDh9bqsoCN0rW3xztQOIXX276EoUvY5h1PhyAyFp9gHD6Cb
sprQaQhl0pNg9v5IP8Bp1ZU74Z6xb2GSAisEEbNzEgvZYDwC/ubWiLqEI58ipVajlwnKBAOpgLmD
z7T5EUYoOjy+rh4iXn4sFG+ZPfoylEPqYHhDWFoV6OjGpgphZNXvk+kwtG1KrxEwcyTDW/6WH+rX
DnnKgB7io7gVlOJxLu+MSyi2Eu+Eee/XoT6dSMCvb9Hx3MAVo3EZnF235j7wrcIyxewn73bzlbjv
BaeSjWlAcyvISIvjxMLemUQBWDR1YIn+rARIu/lZ5pH+RBOhoTatMNPBcjPHMt2JnNpR4ALuW4qO
0r5QDu5gSYZTGI0le2Mj9sxDcYNvqNsWG5lGvPkqplbvl9nxX1r1f01q6dIbfg7lfHGLHRTOmsi8
gVamS5iB2fOnROxVPvcl9W+RquqHJ+BTxmsVRwF1fFCLXq7Da4+e5hVc2ZyAIfN9yUxA+GnHUgd+
Iyu8nCJMmp9fgsHWTI2fFt2+4PBLRoQxbVtIO/0UpJuvPsK3bC2qi81jG3lSjh2RQr4UjLJrWoMB
qolIs/XkTihFilGbj2edkdK3NC85veX4HbNbJT6i0glMf/csZm5WiFCT7OglVHGgjXMsCDRuReq4
bsITEYgE/3Be4NxZtf8F5+2NTpNLTtcKPRO5U5XUw+DtTQQsh/kKtc5zFBQHmy4OFDl+d4/Vgnpf
Px98LpINamUlWlvVkZnI0MCt6f1MCMEiDKUBT/5kzBhd1gGHm2Ezq5s8mwdGzNvzsYDZ6ZITlAYg
35gwlSlqPj9mG63OlQZfZt8JxNCd6AnKOYs1neGvq1kHKbG//auVYLPJ7nhTSr8djHgECt2tUfyz
pVnqLoNlXVKKDn5bnnMwuCPBcHVIliuAq7S0kIW9qOSoNWugcQ6H7wZU5xGpVIEuw3I5UUb06tk+
B8KAfzlYacOKjpLpQquYiOVJ2co5xlJZwqx3PHn+7qLcIDxDRvsgaxpeDsqMzrPy/u9MnSBxLDXC
xwKkz6PBP1n1IDhx53Xn1s8/1dKwNYAe4Z0CXLxgamXSjrNWXpbJ95FRffm7XwjC5DCzKnrq/jSM
SBJyAiwRYMHoQ9zkxYxWGv4bqj4d+V0WqpGzu2crgFryBpPJGOlF9+0nSakJLKy7BHIhSiBAeBGq
yEmReOy2rFVFCfUZZaS4bxaSgg6K8ftYM1VzlcFv3TR3vG7qO3DWLPvaVlzdmJy+Wd8PATGGHGt2
02Otuq4JPtfoEDN//c77ocXLmM85ppUf24BcUPzTjOc8ZsE1BXxi2/M+V/aDmXWkVP2WmdhQtZNt
u0Tb09eCh0zbgu+sWLbeR/Xb8A/m3kxMWjD7zdl5fe4W3BKO4rf46wiocg+PIC8p1aQCJW2HVk+8
PltIrVau1pIAD5GhFM4pf0Dm3Eg1FHkOROnt/jzj97McIDAT5GPI5jhJbnItrFzm4XAmPimM7EfG
fDSIt06nXFrMHRFoUzmhU4Ek536TZ/GBMp/nvVP6DkIJjEQ4HfKokqAJVxKPfegOpWOeVT4wn93v
tCpyZBROexvh6j3TMsrenh7+G5gH5tYr17iQ/S72sjteyvZ9MWPDe87VULpPLMFGUatieHm75fWO
Q8Xmhv19QNO9Pi95v5gOpAFXnghZKy4O1Dg6Z7St/4bUj7PPmqn5hLlr1Ou2qEr8CLuK2uDTAwf5
V/aDBFiYw0N+1egj2Hhp+CxSxKHFzd6eZEUk1VlVA9p9UaY1R69PjcuVdnxRAyvSds31yLysI/VD
WViZ++rdjQIwL3A03d6JSpimpSM8O3D5Ch2sZpnIh7IH3PNJv0mQjxtdWnNMQjO4NaScWVg+PGOH
Q47rY59kUjXkA0+8xnRx3XKZ7GYCcY1VyCqhvPqeLr6QVOfkK8aCoPvLARzZ1MhJcM57qFgiVo0g
/y2qspL8S0n45+bgifnAf49RK7lULKdyATO3ocF0SxMDi4znwkOCOdkSu6FdUcmbLOkFO6TYFpCA
v0FRpnM3vbMcaMljSW/3R9mVnoD5bibRNYy4ieM+4KKSu5Oc20bCZRt33PiVCL8f7vquPGY+FyTf
nlroQUBu9TsOWyixgGWaELunqPBDNwO65yd3YHv6pvwRD1PBEMqR/uwcxAgevTMCjE+kcMGAXukJ
LAoNXzMAp1+MMdLRYvkWinznWaAUuLur7Fe5rrEajdrYku6SbKHPvgda1OYtLlZhYTJTachALJZ/
wIL1/wLNTOGQhUpapF4NPAwHo7O2OcIjqDUUq9qu374dPP8AE10U/XFcZQSvJC4oBc8oZsO32WfQ
WEFdDDc74M/OfRNocXaUqUbbud2ZuA0pYbsVZ/yArsb9tB0ZUTslSGt+2JEIB3FR8ZRPy6CctFeA
9fYNSV8stfLaWQpFduYcEQ1JbxWlqsHcel20Czd2RCLhp0CppHPC1Inrv5+xh0hEjL+tbfyKP1oV
sLPB5JIxKA/AiQWplP0A49GGOD+VjCi48oB1EAQYlwmT93mrDRgwXHXlNEC3S/O4OUgkKxU73UOJ
PRsmuGgj061EaJySNOVtIZhPgiiknWtEmTvkOBgk/pyXFLs/DwmjjK+YAEe6xC9ndHIOva2fIAs7
xdl+Dia183VGSK4Uy+guUUMVTbM+734gTzdi84F+s3N0+928uX3QTiTUhoJ4W5SNuFilB0WUkaEx
Unmhy26Zdz7mQOFCW4dsdqteMbYP/fnSBEGEPt2ofUIrwXd/ggaowlzkPH+c018mebSVqEi6WTbB
U70/8WSaqEswVyHbkX5r4pSD+YYMEk+VNVuy8ZfmwZzu85jo9tRPNurq9m35dsZX/N6CFCTD+lto
cHlcXI8X6Nt7eDnD6qMGfCOYVRG8sZO/ONSvEDRGUi1xnl2knZZ3eKRZMAmNAy88KSL86wCzySFo
22JWQzT0TPnaxD/N127VVAwNcRaMSH7/T9CB2dRXxuvMq6KIpG95CpSsUqqqpOiOH/kiEvYWliIy
y75FxHYKLoihLSgyf6A0q5CapiiJWQ3d455H9IscAVeb+/mK52naiRmTMJmxBnmNXSPM7hIAk3FO
1ilB+/IvUHf81JzOPfxRi7dqGQBz7eH8l5ri+SR4hZpuaSra7aHhcBauXS/D1NpVPyYcBvqgMwZ0
BG+C+7I2hbctp62uQMc07XLrJfPGWG0MkJ9uqQ5yEkUFjHYInGpfkkmhbIn7nqiELA8DLrU00cTY
586RKYrADGKxGZJ1ybqyeu5igeYAABCwI6++bGqjUr7FI87XfDCl223/+T20xG/iGS4UjPmeQcHH
0+aLNxtU4AfGAneP6+pXqy4jwACE0lpcrlCCHcvcJRJwk/LzvE+e/I+pertMBC9s0ag+j6wopUM+
hUzvWbYwmWp45Uu3bS4QW/d+KiID7XTkSkCQAEdvE1rUBKVwhsC6A3kT0we1NF9rG+3NjFjHHCG7
ex8HwxlQE6Dj4Hra/VzjNZVe8EZdKwAKbKghLCe4SqqZAFlGnb3RPw5uvk76QaWmDu0aU3E2CQFE
THFxO4/K+vx7UCG6DZ1y/KvKZ73HpS2W1LGUPRuABywCp0HzGkmPYSkv5nFJQCgz8omi4FeQ1XDz
FKCo0BpcUDk05mnwzgFFU6jSXCzd7JFd1+FE2KOuRCV94btcz5BsCUbxd/PVqH/CWLPew4x0OxEk
8+8nN3bjv/WNaABmjvOCJPpSQsVoCRoEtK84TbhYM1oZvMvy9IYzfN6Xy4jdSXSpl1TcZdCgXOkO
pNS8BsKbxo2XHY34q8h93M298tKIZoyAtnoLkK1qHGSlhbDhhF2fSMSsxPiPig47dMTjOUP+Etrn
WzO0aTq6T959GofWK4TaiJ/0yXJn+0AEfagH92MnbL8w2tZ8kMANmYu/Wn0HAd4DSWW1pNZer4cb
rCRqn4aergMR5i11XJfAyyRJDFSAD5/OIROBf/wHiCZUoc/JcLSMadTxW4US9aL9HaPXrT0ERFHS
+CFieBimTG0jJ8LnfrCeqfO5vXv6LHaEOdd9x1gyHpj+4BG+le2664Gy6q3jgvDM10teUgqvtXO4
/friSUHlekJQA8L4FBUAfpeokuSgPxEkTiV3KgfzuzEApZbuk0Tb64PAHvUIqOmiMICiWlk9cbYX
OgtlAw1VYURKmEsE+mkePqU2O4i3b2GhMopqivwehw5sCnhE3M+bDPrimPeTTevQ+73zAmAcQi58
32nBvJeNq9/dzSKRDqRMPAYJ5Mw/cLSCzx60G97a0x+coMTxJSp5zDoqgj7xbNoW8jNtXAyUvhlB
mKWQC3R7hCX94Lf61JnMTHHIHJJBucLPOqIbobE2iZnthsOR59wVnmLsXx8PVevgtpjIDmcNJUBZ
WoUw30Hs4T0h7pwsenzz/GHDVl2UzGLOZKUdjwWLoIJKUY6LOk+ptOaYNA6GPqd0/9GClmKoXxCz
4QYtIUAwHxTZe1ijDm2HKsaPUwoL/ByarA3gUB6FxrGxZQWIeX7fUvdj5cOTnK0weZDLrjTTzPK3
bb8vy/J3hqFfRBf42mqsBKYZ91QXzGRs4JyvP3f6KYKwa+SaNe7LbO6XOd8eJQBXBicHnspfTye4
3J+btYuTOF0S0NUKSOBfKex2RPGQhFaqyL4mzG9kcK/3Ym4fJTI7OUbKKJgYlp+RvJATdQHjAtxN
1kZtkCRzWJIrEJvYcQsfZJo09yy84XH4sG6clWD9NJc0Z21rHL+kW04TKkdpL7haVlxE+imqmKtV
u50uQWTWAKL79fMmPTAyVA/IoJBHB90W14VozgYx7XFzDjmkJyGqDlcsHxbLF2Vi5WVq1EKqC0ai
71TvWTuWB4oOrJGDDvoOUy3TY/Czb7fMRjnwwfMyrWi3HvkUIH0isdrO5CenC34HQpvRKhRAm/hX
wTpvcgoDMhIYmSBP6ckZzGMoJqcGYt0no8fyPKaGEBTP+bvHztHzpmAk750AtU3MbHdJKTXk/ESZ
75REmT0RzesaL5c53SMk8yYXsJQdMNZoJOBgyJT6wBerRGd9vMojwN6VMhMRsrmJSYaLY9TwmGk5
/CNcXlM3M3KKowulTZPQxrBjPH2Uf9wPGJ2BLasvRlido0FphH6gcijxEc+6Mc6oNgrFEZXy+E0z
6fJuL/tR4U+amPPASCFqkeupcoLGCuQDY4aydeSKb9JJ2ILo5Vl/iEpxxqu3nHdm0t/rXzqwEt1a
Ptec0mq5PhEM5086yeMBlmsNCYt9JJq+qtyEqOgc3fTjZcvWiZdrcO1ZjYX4E/Nr7vLfXJ6xNbEe
Hl5iXlBLIBnY0nRU2WyrzfuOoIpNXa11XuX5HqZeiGdbp2z22zB21w9RuFuTcrErUq6aVkjEMvyw
BUnTwdqp2P4VbQxeEODX2PjIaXDAtMECAP4j1nc2Z0wPoquekAURF4e02uTMcc4d5xi6LbMaUOju
CKsGBgqgNzt47qXoYyhqE2Se0kTmzIWGsBZA1qNJzXRsoseonxqk7NbwO/wl7/VjZh2yP2r5/mN3
7Zi5nVhpDDWrG+lvpVkhAzmE2ktcjQ1LweehoYDLE7QpyzAW/UxndIaTh9QwrA4ynlU3Y4t7orAw
AwZIISypN9IyFPKb56lBzzFmTmfG5wqhfYkfd3a9suYE5o64Kd9QHOf8qlMfu1kBpHChPsHyhuPi
iejNosq7PHb4I82vNfpKJ4izcBqGjavm9+DFPZc9aFWN5KBIDoAHcf025+Pvzx2P8+/c436p9BsZ
MMpNbdu8zuWvewEXHEljfT0fefq3iyb+NeoqZjeG9gM3feNRHfj3gibitz3MilHU/KO0j+BnmBdG
EQfD8Rj1Vfg89IPxez2d5Mypx9kWakDYDpMI/cHAOx2ELekuBZFOqk5VY1TrreiorEzm6eCBPM4X
dmdzJ/ubvJkSEBegB4vxTPayjS5XDm/gZuXjUHiz6Cfs2hRakNPTt1xINF9xbtBymAlDeHpdY+Ja
k/mAmlsUpvtZaEU/WkKgta22yKnDcT9Hid0kTqrRV+MW65uGZ+mdfMArbGZ/xPiYouiF4/hJvgpt
/N8kmjm8EbGWuJf5tJLkR2CtqYA0fUulcco23BDOnSnC1se7i3y0n/u8JJT95m4jMgnIaUIMPl1X
wV2aOS5ppQ0BynF3Ha+ROhiZ5YR1phaYLsXHIxKH6Ka/WP/a2b8TK4r0IUDw8EN/jMTvdA2dkrwJ
G/mYgcSL6qcZ0gOE/0U/AoiNrsdYRF9DyMj9h93osNoaS6dQO20kqQ4EGp3SB/+gtHIr+opkbVyD
NJnihgzFoxfD0ADxdK7PSfWA4G98lOX3lg+YyWJ6z9HMZYZcgozZHVTSWSZOz5ZqiIh3wExwVVOo
zdviQ/awy9a9VXsIjFy8QKfTjVPVx+VPf/93B/Io8SyHZHDrtlgrsHvee9GDlXFvH8Q67GNDUWZD
78pT1J+shU+io2mYza0DShEvql3tZW54aH5pKB3IDAUxC/SoFTgmZiB7j0VY4U4I+8l7gWj/8iev
mYt+6hUqjpclRzxsR+XXcGYERYFV/Kh7LfWMG7Q44tKZaSIv/jNMyqAu9BbhabBqsf73pdeLd9ip
fmcepw9yKmGefO0ohyjAd1x7BacxCeuaqc+c2wFiqYRGV1FBHZebYZfJPLRscoouoqBnwgvYKUV+
N5tCoeF+NIdje8vpNwUPIQJG1ysWzBjHstO9XggGqmle2/EpusFZDv87EFezS59Sut7CWwERe7+s
MiRlvneziuq2ENn0ReCy7yU+JFkWmsCMCAuo6W2Zb97akrf3rNwP4vyWUJOivB2aISZwZ9/AuM0l
96s/VuyGejBfKsu9nTiD7n1tMNvmg/SiQS92ElmlWFEsT69Y9E5Xu9QMQShtq2IOxfBrYQ1lQOIm
Q6wr2cDXUB4QfIfHfenqBa9sbfWGGCEnUWIl7qNpLoWkc8BNzG4rwQtNszC91QsUmVxe6btoqMqv
IO6dT2ZSIBK1F1nxFRK45ccAX078RI3eFxuASJfz+d7tDdVw81ffDFX+DJF00E8ep7uQSvDFOBbA
XLrI9tu3y/GYXDEUHTcxYUHwMwcA3eIw/zY26ZVRkpK7HZxt457eG/sff8af9lXMhbKftibV48fR
Mdp3Cq6Co3kNwIAXIp/jbK2gIszRPphdf2UwFlS7P+b7m5+IlLobUKNk5bvPgd7aAaHSnYrz8b6J
Bh68ett2HSCT+7IH77NCd2Y+2lEzOofAtUr1Smg9CDuXrqqB+fFN2H2XcNrvE2vt//bYOn9JGAn5
Li3wA+z17Ww7iQ9V03ORjVj0Gnl0vZVFu/CQ1TP9LgYsjV4iscPqdP1rVjis9Qw4kYhl5DwJ8QHP
koxi4GVo5AL2BpxkXMa8UHmQhCySbVsQdRJlZrtF5QJprwqvYTwTlQtV/t3KOQdpYKlgSxWCYa7f
+Dd6vN0EYH9QcbsDuO0eyDxwg7+NoJKjuCNVTjXCazeFi+PWoSdZAf2B6lt4qU0AGLAFHH+T88NC
LplBj/BoQzL9V3pMYdxXg632BYlr07Tn9XM6fVkC+xE6uwgfJKR0H1Tvlc9yd5vuImEaM1EHqRLo
Ufi99iSNJleSd98tS6+rGVB7Y3D0lFAkRhnu7VTgzrVaA1Fgif0vuUicckqSTWEMMBfJw6wEXxF5
JCs4oIfGiWP1zkV0vNklCKzP2LCUHYfHuYwqe5mey59Ye/+ALvZVDeYJsl2We83J8DWHPJH5kb48
osS3B2cULcRkSFueiYdBil1TNOXfQPLxqOmsHqYkuZn9vqhxpdV4QGtbF/i24nyAoyyeHcBHEgyR
XOuHaYKOEgQOi6TQclZHH8zDG59ZT0MYM/HFnUELDMYjmqRl1RnKJE9/YnC8yCZ9a59/Yv9olvPz
ra3ZU0uZBTexjenPm88SjHkvZOytSI7qqt3MOeasVhJFZt08pMgBt0bVj+J+r3Mepfm3C+iO8Lrk
NqJ2Cw+l1GX52k553ufQ4WNcfff4nogrhNEhdMhbRG8f2Ae+xiXXRCBkrAVHNPnXst5/XA2lb5zF
TRY+uSjfKR8gawEquk6OIi9huzZOm++5OxWcF4emL3hb3Gk1nnFA7bNOG18St2dWpQBbiYB25jT1
43kcYb0uJdq3e7igQJdat8Z8qCgj63+hDJUn6cIhHYyq1mAAMaR9GrSAD8A+erPTW+m/qNpuhpe3
MzuMvEtTuvdYw33fQAeczkmGhWCOZy4nFNDM5I20hUVw1wf3PujiuzKLs7yQLSf+5Tohm7MAYPIB
Un1HcHpmLaE8KaJiJ4urYZpbLKKenATv67JRjKhunK+bb4OgwjpbBMHvsHHrrChjJlW2KXDGPnAl
LKoZX2N4us2CXhTJFquw3D46Pwz5Te34WWXgxIOB8je8QdKe7G2ZtcbNPn4Z3MQQx/3/4aQynEN+
qhcfp6XiRPYyzgojLTlzD7m+C4jkpZoIpCy4guXs2tmL6MeRVfoni8U+QRqL2kf7Jm6lxdCMz5LZ
jn+3J8kySrDMsz8CpGWmXy2PjVVx9vYdKSZ9fhi3/k24bpaKjlTMuh34TFevCOKIukD/uFBFZHRB
KruxcEoaIrXD0e3cKyKCwhB8m4fxoCirCk4RLSEeWo1KTNqdsnDetCKHJKxNpzxaUlSBB8knjlFw
PpHyk2abppa9IxhdRQC+komnyywZcZyHYpDicrjVaiUlZoTvHTcWHWt2SJgWXekHxZ/Z9fZ+3gJJ
zhT1FVxx/fEC92UKWfukgU9qF55P0VVtfc0cP0M/KOUG6pHNg1DdKNsr1wX4+Xo+go2IydnZCs7N
iCRh6CE1zCYr8u9P3iPaZqecK3Br4AGv5q0Wtl9cYxKNjvUT4D6vMKmwePEEp+ijE5INNogC+9Zc
RTGNJJUNCTvVQkjgme6KhbX7yv9EGdy6auz8lm5v8pqw1Cts0hE2JAqsoZEtnsPonVibeJ/qFneh
kzxVg6b+Et/syDfmH1sSPw7BA5XoLbkrX+ZMIKQeBCWzqS7IwW7RTuhh/y/kGzBuFfPYF2+qWs/D
MCRXoJdBZKjlb9O4iRaU6MbzZN9NAeBmcqBvaNG2yHss+1v8VZafJR5hZdv21CsHq8D0HvJ2gwyA
ykZ6IkvWeRs2udQ44CN8LRieHTWnnWqQ/8jMYtkbWEJSHH+KcG+4r7jxINLS8hDufNOGcKdWfuxt
D8gI/C5VzxZX7K7uUSDZ8Lh+7sMBxYCOBAW06R8wao36+F8nOPdukQVh+LjHhN5jNV04ONH+2NsD
i7ZmUdk1a/Zj+vyWWqBlkCQwoUYNjCVjFFfwQNltZ1uoOJSqFBt5sbBghfOEBdDg6EUaN9o5L144
mQwBYYGxoi8ZAC4o+xC90t+sdXV/AVGcBcf+vNg6lSeGt1wIZ5RpOxYBCEsLNsKUwemhiPIHMN6D
MQSZBP1bppH9GRqtCO6bEPMLqhP96iHrc06q8usKrW2MtcmI8pM0oYVfOqJpn4NbifZiIgFWWEc2
wkjXE8mEoa05hWJYITqwa73/yRKBITgHGGVcHvKqUY/UN8ywhhqQi9I5lzbiXnhOaf/kNdZUAUYv
c5O5eE9Dr4hVhiGAQGpOjKHcuvxu0RhCouWt0bS4LUL2m0oSshxXUbH64oum2NU5lt1zTQnT8c6B
HKEIXwAr95n37u7xE78HyZvpbGjaS7Bkc010aNP9kZNktOunYOL3NAf8Ekp/m7LLtpR30k2Pyy+x
el7XID5lzbLveZ9ghWxsc+BbN2A5M0dusJCskJVm/5EvUtR+/YjzX+jmCzZ1MR/tGhhy159blwjm
8o2zxsVyTRKF/+vRkrHVbUsELn/SG7b0fzs9UUaY7LQMAsEBxHLkLQFp9iZ1H9a9lCYQT0a6VF2B
5PAQ8YOOsgqr5pOXF3efoDtfy9mfqmCsPY6n75XLhcafooTouupMrx8uSWT4kmoiViawSonJNWKI
Pku6CkQ967ODQ3/0V2dYE64JRhcZu9YWDNYmWxhuQH5hG+cujiJtMu4SheLH9r1yoT88Xi9OhOpS
+tJQCdxUIBVeFbkGdX4GTohFRVs8KnJgpWX371b/zAeFpRGxUUusgH7HWSbQX9H7Y3S9sGdLpuAr
aIi3FOjG9orUHjJVvooQOsReURnf74Mks1ctRRF2Ea5SFviDjiq5ZqR8vl7TJkNK89xQ/8ROoap1
ohz1ePNQjR0QImuXTrRdPtP8jMS1pO84D6PndTDOwyQWC2MDu+Eb5ygKsDq4kKQoNE1ka0h61HJI
C4/RrURSRVnxzo8uff/piGWnStMVAd18qMBPfSdEkJOZBbBH8KU8O6l7Cv1DPE7dZF+QsXAfOpuj
1E8p/EYTSpGWNe0r6dtX+602DZBfPvC4nu/uFzoTEUvtTT4S4qNyA+pk2bYUfJ61s5/jsjIqkeI9
jfg6zy1KewsJWFF5uptFl3T1x68BsCJsBY0qiDjPdf8/0zJRefNJ192aq2qKxqZ7bhj2iwe1FhhE
4w/TlO6Juc7wS0J7VUN/U1sInxUgJLNdaU7f1+YV7eXrmoiI/Wp5ZyCPERPzA8mdaTBaybq8RDkw
zARCMoalXjWljFCow3g9qofVbucT7S0IM3WZ6dPgDAlxDvW4gPsEQ5g8VwLpqkSv08jbLzR12ji/
0cBVtsrs5g/V1PC8o8j+91sjXZfjp+qoOmKCN/sqK+KboBFPIBJKFMXQu+LV6oatx1gUB5ujttjR
uqCWh2Wr0vbAji0GqMf60COevHoc2IvqMZ2VL22VLqcW1FS9Zak0hHEKeglBGBqjADUcJ18zK/HU
brcRcqf1XoTal92JgNFQZajzY5s5B8AJJ45UDqQ5fqnLGD8u+ZeD/gX2jXNQe3mv0Uay8ueiEfZh
3i3EXtiaeVdsqpyB9l4sZ/tXnrbBjVKgqDCxOYyAhB/Wm/FCk3AaqLSCGB9jchDrnmzvOQYj+xSF
EN5yMYHUvLzqro6cm6hIefCpVOmKDP+x2zj6fzWlf/OVf9l+Fogiq7y/zPGewtqFePvPMS5l73mC
rkWrfBLVkFA/QUEYN6CN7hXmP4sG8kZFA/5gs2nHGzrF0iEMtijjc8CcXNQ3WBoxZ12j96j/swn9
vLqafby8JEElBwwKI/++0cujikO1Mnnl1IqbKOA/CPkdF2tD3JDKXkGXg3qrpixA8pTm5jSg3sBx
e2R4yzEWslkpKGvAMGZEk9IcgqVsoDbOYQT5uPiWFv/VBogyGclff8WyBycZYOg/Pg6QyDQwF6iW
yIYR5AOjKBcUsCyarPFT1FCkylBv49VG4unWUl3yBC+bMCHdbZzh/FprsqavlZ8Vx2Ikf1GQDtTF
TgdBUdwoqlTZZfXJDdB0qMisucocDBXerwlTMGKtp+fVKOf7G8Gsm8wi7PIhZ0rWjiMcUkmJrTg+
mL9ZnQ6MWDvwBhurMg91kPF7SCsjsXJp3IwcCRllH8IzmTZnaGz7J+UiFBUBUhVpm4qKqsXIFWtc
BFY+QrVfo7Fu5dv61YQxeqzei6LWqOEw20UIcUac1VFkHl6OHY0QR4S68JYOR99CGF1z4EFp7kwt
GxHKULWQlKXnYz5pOvOG1RBdh87dOL7ln+8vAa0JtDJUTlX8aDhdJDIF/BjImCPSEnL45bdXU4gt
udnkVWemuQ4I0eWvOK4zn5MlveGZk1uDv4hRawl31pQwQI5v4eGV1rCE70Xwo8nyViC53YG10iSc
HivWszvmyOuLTtXCOxdWv7qDRGMm7YGseO1c2Ewr1MGjaTwmO54JQx0dR1KuWDulNoQIZCKoFY/Y
fjHp6dOA1maS3ikHkWVSMN6oABT8A2xXrkp4vt3z4Q08i+ipQHdbA02QA/7aBpGwCRIsQAZY83mB
mg4mj8O1UmAeo7TriH3s/ShjwiTG7UqoEV09Cfx8jA3kxpHjbc8HD7gVpkVe0RRTQy1Aud/KsOJr
h8cNmuC86OvasRFKWf0dRPjHLMfkfvB37VWn/AA7zTdzXUZTEK5lMfpZ4EXChmsAGJlg/KatcFbJ
/KBqMzkm6gr0coE4jahisNyqXp66ZGkPwNpZOZft1JW1t0CBrYMPLYgcwgqtQL8PPAmDzYf0MeBo
a5iYw4l3IWvtn3CMoh4arbAY2AMHQBQ8pGFSQVPp6Bsjd3XtuC/GQ/j+zw7BUnbrmRXUIDFc+DjA
57xxniryV0KTFbeX5LNn9OtRRUTgilVoC3vbCTOjEiI9uTOYLRzWfUU/IKXHl22IofsQ1ZOMrvBQ
vhEp+KW/maZb/Lt0fgPTfb52TxhrW96hoKBRZ9hKLaK84QJKzn0F+Fs9SG7FyhJXIpMM9L13R4D0
cmUf/BvHFOTuLtaHz2I3YIGJi/pSe4X8jO+PL0NpcDwdJfcn2oT6Ki8osEfVxUkDKb5wspJ2TJ06
78FRzM43h13lybcecZVs+49YgtG+H9qgfIGbvg2IKt1kJ7FOh0iwfK1uDFVIyAHpQwK/gi2j1e2h
HBDhUpKJMApjO1Fdql5RW1MnqTbe5iRAx6dSNCwEROudThEch8VKpT2iMgwM6znATlCD9kEnQSDj
FpELJ0mZhYICCicT8pGyQKH8A9PwiDe4xfHg5TUCX/+uiGLw9xnB80Vct0NIsp97KQbRMCfK0DvB
cfznJferZPjnPnmFtNRDi3dAzjsKfQipARjzF9yu3yr8cAA53IVT6Mwl1vNdXV9AvDRJn8N3XwFK
GOtTkU7xahACkgk6WpKqDShfQj9RjM35M5rBFztOuGF/HtTWDZ6P4yOi2y6Ii57BQwcxvNwPYqwM
7QVPQahlTmSamKDYQXWQMmHje8mrAiPpcbQabChBRomUCjGD1nY5GlrFHDs1lxKhi9FDUtvyEll6
G+I8BUe8fUg165XBcSUkNHzcEdPmMb0ztfFXT+MDtc3RAs8kd5TKoYLzDRhG4NdBC7oOnab8zSJ9
efZlCYef78l8TMmDnSNguc8Fon9WJYt20Ps6F485SfFW/gyvBHU9RDkvhsxdr6hhS/m5TBufw31H
P8a5//uKs8W4PDs1QoXNu/GuPxqq0Tso8xPM9ES1diw+etbzBgp+8qL4HBgS3SAN66ZOzkwsQ37d
iWwHX8JaWvDQFfminsB+MRX1cLYTDwAp/ov3WIm9kb/JuoW6VqeARxnA8jursXVadIgMYWuHE1J8
KAlugcDsC+Lszt6HnB8kanSGcnB1Jo043e9G2VWXzRke3msGjvp2lWgg8hDhVTnZV7lDxGSSu1z4
qqYDkVLWX/CHjtPnbAL6QIC0Kg28q80/lmbxvLJj59MB46zks1KoZlgB0/GZ5lgWSZe1M2Ys1AES
S2yvbicko3Oo/3qvKY6UUJfvhCP8+dIECCqgI2dAPOsdN9Pj6WcQTu7Aw1QFE5s0uTTKUjiyQ7El
6zPLZ9EsRpFptC0UZLP+e1PL4HrF1JSORx0Jnh8xUkgSLzW2iweSnfxMiYTGY+/5ygTF5G0gvV4T
ko4Hvqt/fDVF0pOZ5wvaO4IDREIgYzcQ7TMLYdU6lGSjPUfBJV6h+f7thkzcZn9zc6GwGKR/oTnR
+HpnNLKtOWDXBXhDHXBiUcPtTSRdHwmJkgnYU4UJqeB7yNJ8xynPw/P1NV0WMD69ULT8IrIYWq+t
jSvBnoS61PlFzK+aTF3/dDK/4OU3kruWchjDkTSz7WT/QU3XgPPtzDYMQYr/DRxeJqK2qSFdgWcD
RTHakf4brpMHJRqn5ezH6BsCPeA7DxjEsHVD54YwaiQhafp3BKPQ8Y9F5khBQreew6kZLCbqqRem
YF3u8AjzEKlfNILVDW/sCfyuXzVNwEpbfiMhfCLNN7ziQZnI36ATEnMqMQoUp5XXTD8YA9EvvuBf
Govpnguh0RwnewxxptPDUXEQvUfJ9WgSUR/0k/WC2FG6psf1ejzb1fHPHIr1jdFTMw/u9AeKcwgX
kxPpHaebwhkWVsIn/+CoislmWH+XNiiMW8wH853kL4tIMLKEAklj7FkF++LvWuXBavD+qSDr54yO
w+8d3aAisp1CLnb5CAJ5kRz59HN7d331Hm+H/er+pajzvDWf9VaohEPZih7276AVtN92d3h/GjUk
0/bHNA1pblyTzO4IBnjkL7PkKq86Nz+dP+lHUVaUSBMUdfP+alrAxEGfkONX7RJOm/k3QcA5L/0h
CFj7A6j9AAzY7AgfsAFx6u+PTg4YlSeKTAHcSoRClUAN5YTC7S1BJNHIfx/DrghETvP/GoOqZyU+
wAb5+JL90snoMjuUJ2Hy+E/GNf1l+fYe+OLYUGNYCnJXqCnN/c/MgcSFcv85yrwsDljwlc6MpE+v
kmGtfC+fmw/jNhWIwUGWY3z0CfazByC69fa904FtKBYl+M9mO7Vslw0bAsUe3Zq4IDPW9y7TXScT
8KIvolz47FJpnGkA0LQyLI4K73Vx9Dcfms5MMWaUDZH713Op/+VDYs50a1HKfmdu19sYTSmOIi7v
tMT1hS1sfhSEvDejCYFvPo4ex7aZ52lHvk7SHHvCxLu69JyoDy6sj6eXV0oQAEmcKeRbbggQyG5n
YBDoSygWhn6C1T4etmRKtTpb1lStImDddbFwCSZgszjF9SXRl0JXJjCKEoy2XCXuZ4u4CmUnTsxQ
gWosnZNcb1S9hp2ciF1F7Sh0qO3YKtYcjBDqvqmh6XL5ptTWXHILPiV9TUnJZg6LEUzTbv/MsVOi
adpVa8JFeRp7tQGh5alUa5uX+571sf/P20BFPj3n8PGP4xPc+gL8dM1pQOdbqtKh3IUUOucEwaYN
A6rg+zabjyQSDzK9Q0QamP4aidkd6it8IMuLCDDVQmwToCDTSWgxWcJT/53rHBJkY+nOgKz1oDQQ
PlCx0aYZAHZYMvZra5k4IMEHCsHmR56iD7+BATzGNcTpdKKmEEErVxvzrgt/qJohykJD7rINEacX
7mMkNaAB0+L+88mVDiLyoc6IqBJ7lEo7xndmvCWLnw/Ix2BgpQ08IKDiIihoK8kkZRDgRTQNXRBK
ynGdGlAu8wPIpoQq+bVYjqFSVg1lzwe0/unAm1uGTGv9OatFpSYRh5i7JV1JShlKhNv9+CGtj0Vt
k7jusDdHCFjxlicsuyF8ThVvi9WaVox15y2igX+HB06BB3ghi3Qh/GJTSJQYIWJFlVQucT+fA88v
Ud1Sx5Ib7gdwLm3oTDhvd0r4IuB6ne8BG8w7FjKVZTd+njdPNGZu9AeZRc7rMRVZtS6r1Q9VHLMp
eIuJLW6TorV4eh5Lt0up8rWlGs0YY0fgVbV0WZLFB7H6z8ghW0RZbFUKnwANwHFvF3h7z7ZTKLoN
UDH/zxfWhblzLhEz7c2hCBN0sjHzsMJOUSh7xOAIyJlg1ZcBGxyZD1KlqfLdkW0SGr85Ja1ueY3I
N8GWzkSv/j/r/IQToMHuaz6zPEA4sEmWRRK0L8DK39qifFFK7xr9jWgbRDCewxcssJp6oPs73Onv
XgPT/2bcW7MSandxTYLEjRWgYuWgDk8rHHLDhuiwVovKZ26bY9oOrh/kcJNAgdjJ82wyZCZI3XPB
u4bsV8fMRvgamhRZ64Y1pQ3GGex5q2j+fxF5x+4d3+Ch9OOtgG+9GjS47/QHg6vbhN7aLYqII+O8
2REE2Pty9nhUR/RgONlNK5qLyxC5BqSTqqCabDjnWwExuJMXiIhxHtoZ/x5quKedhoUl0schzQNx
uFrR68DQ0OJ9XABNtL2pGU1gr6sM+F4iQWFwwr7ZcZZYmxHpnbtke92eEXVTJ/ifL+DpJnZD1Fmh
m+sZ2B6hVRbjKj5+2Rn7V38X8lnw/MuCTC15QRz34H1TCnq0BvmMO0Cw7l8IQIIWbbJQ5C3AJDUd
3uJuiu8c/UWnamfegFU+bou24wbgACA/joS4MiTw0qdppmD4FrtdWmc06iw/UNVsf2xPPyep526V
bEK09v12JQGpFle5GgeIuEYhA15yXgFWcykZ3bxjxe6jNCfxI0cyt1roT4xTscIVOmIE8IyZ3uZN
AM1e67w9DO3TSAsQ9HeAa4yZ/w5mVbt3brvZh5kbOa7QCPI8mfocYoKDR5yEctnW6DnyM87u+GOv
BShmhBpTismuiGETgI6nWy8t4IE4ZliFJmB4B34MkufLhGWX1isKeft0oDGIuKSmpanqlvLRvcgn
ft7uOkQ/Lzjpnlcf9kxw5bZzNh+gMODPShNP3KdE4SY4BeRxWAvXhvCcR4mFll3Qhb+lQuspSnJj
Wi4djPtEmiegPCpnoXuI1L5wg2+dkx0Ia53FI6MFcu+75Z7+AyqkD/iXgn4S27HTQ/MVrGXTotNi
kU4NZz2uZlgbXmdyw51B5xD20n9IcZmqlhUmO5oyFKxooS7t2ZvAP6Dk/KV9m92GZBJHuxjIX3Wf
iLVBxxTTJMTmN9I0Asr9ZcRZ6jMoYrwE3OXIbWfKcv2xF6NBELo1s2+e2MKA5QYa+ftQt4Rkvjlt
wPWDGc4ZtKxmNZLJ2yDZd518KMKHTmvkPkpADEe1w1TgzQN8a7kEZdNEC/S+xQ297yLud493oskB
gAyFEfak5UYrWnQkuFwZBMhpi98YW/UIStGO+PcmgvMrwPXPQjvBC/8R2TiIjt+UnpOT7Ef/pH7g
rXN2h/ziogwV9QJLlH6UDtLIZpxitIpCvQHivDJsEWpBbGYrEq0ktjtm6rW5pN8ry0YybZJcmcDB
+XUUKYrZkecKh9ilXxVegaYVkzrnhGtjTgpHOMuYD4zfPVtuZlsMoTDiQnFY8yZRwQEqnOjI86wR
siVPvNo+3kZhQKiEM+jiRIY4LN8IcSzIb1dT9mNMLOHXjuIc4fABvH0jKL9Ju7VX6sWkjnXT1naD
xMP3ASdqoVjanHI3W4vCIe7MtoZ8PuPk3dGb4GZPjVLwyw4gWk22XFrPr5DUElBF5x6v4Gr6fIZ2
AugJUNbNceNlkJ+QuAHZekGVspsOIPgdBKrgqFMi8wrHNdIThAi0No20SJrQcDVPBpysOPRGjuB4
Tf7+cVjL2rCiZ7T50m/Ooh4jwq207+0NLeWGKax3y6i4OpOMVt8wZ16QrVYWvNsRkOt6a25/wXO2
4K/dCp4KMvW8CkbiMJlXMfI6SCG9V4kS4ocYK9gtnXde2V0HnyQuly8N0KySwsqiswJ7nVylyFZN
hJrQ4KScDnv6FIyi83iHOnQshK/ousfMR1zwhzB123pZosFxj3VkJXn8x0220r6+abzSS3dBixhu
5CgYyBsUEy4jfNJkEScyWwFfrYe1WxiMXYWIUnmTCCB4efbQCCmh5k872J7pLOK66tdb1dV8TciV
o2rcY9Ji1KCVH1CvCh7b2FxWRhT4BmcWq8PmUcmPyEAOx+1rUxkIBnJVxkm4tYdz1BLynHib9fN3
KrXgrLLG6pVobGYGzlJrjET+kT2n2cZiXJvW1t+2N0VvfdH/JBV0v373TsnfwjLiVbpPJwvkWlWS
6l7ojSzdaGlOhsm2aVvdKwogd7DaDfMuwE8rk8Piep/CImCdGVRng0Y7tcLjfd2wBp9wxFTXB6LM
TQkF7UbCVV6CwY58njAI8B/CXyc6L0TmYS6vY9PSGxHrw0nKLiDMHWOCsITlqYPbnfC2u9vb92cD
rpVQvK2bkF5exBr9nRUln49iZL5Phv0KkARx8DTn3HjHQ6JIUHhowXlz6/fP8y5iQddJncvdHXEy
wUg9rMyTFpd2qfy1Es0YcWE48sAT7vfrD7BoHO5wOxxDIwxZlJfeIPOBVXSsBpUHJQWhOXWDZQ0y
pSwybtMc7fmPnCVMVUY6ocZ7GjI7lkrUCVfhGUyqcgrfuHrogYgqq9ddrdB0Zp18CfiLpYS8mIG9
yJTID4lRQKhBCOvPtcTnKQdTPWT/bmLJ9qiU+QoTCSpRq96D19lfwa4UidN6yCnMKYcDHNN9iEBK
kJB24gy2rAuyXXQ9qJfThi4U6/OOmt9cBEHoSN88wkZZJOdsWOw6enSq72SFdokUmd/ZZrsH8nm3
D3HDgHj79DM7a/31DS5svLmfjURD6MGFrt2d2jhtH3ZNtkOAngcFFyDE++7OIGGXTfFGAX8jpk0p
rcuXdC1caF0HCjl05m6AQzg/RMy2+ENPxKFS+F49P4cKPkTL0/GKScPr39rSHh3WvP8ZKQLHs/9R
CYLT6ee7QBbFmJ0XT2TX9+ArfWqtrYwJ0U8Ptc+IAgEmR5gfFlRHEMMFSPb1f9GC8SmDLHLR7rr7
hZUWf2SIGZR4a0NC5DY/N97tQlPfVDjZJ4Tlm5cEpcvOiQJPWQGTLfj8qaUKgAF36eWR0gXotsTi
bM3eyhlz2VDx/E6dLG+mLSEc5W6JWaLUCTBUY4IaNKKVTWTzK5fNZqKGRyxpM3m0lm8gpxRB3GDZ
nQtD1/YKxUmQ6XpFslcNxjKNryDlOEODt5svLf+NHs8qnOpS/ccCFdHODer6H6mMXnTec5ZaUPvS
AXzrlZIbD6m0+iw4MADpMThqAtsjHE+QU/Lx5XXdqW0ZJSMHXHPGK3o7FrqSmGIdSe/mRnQ28EtI
Wn1iGZ9JrkJMl2lvA2ASorWFdH62cjWqt7S+9MfEsBjVs45KbTYfMUbGLiV9AXVxpvzInEIieDBx
WjHPTNlT1jdr+P9/312bZdj+TI5YDDYLYuRt3Yz0AR5R2UVE+kLLgOpMxWw7N49WzwbSLyopWYL2
lJxX7cGRHgKQRlodzT/MfMZ6pIQ8HCN89/jH4ZeYh/fd4wr0O2G/5+DRsKK6AoSejpU1xMo3uAqd
1XyvP0j0KnhsStnPRYuPRBz8uZUx1Z9PfyZ0meIUUGp+SaIxxGYc7yGBOvTYbIUJ6u0Jm+S0+30U
s18QQOkkmMi24x/dTGKxBxNL6jrSi2PUEpVAMwk6u3jWuVgH4XSbrbtImHSPJR5I7tD/XvhXbZIW
6Iaz5tMC3GYnHhI5IiaNumqOHfk7yC9ANBkezSs0L8ROGnfTqKS9cGQYCyy1Ip67YV3LnYdw5z3l
v3Uu5c6DAANMTe4ZKdVdRF/wMwPzsSQLiTeX0BH+FRvlflQ7gvWPRGdYxwsgcE+Aq4mIm50HrKB/
0Emwtian2nN1Hcpzz/NJeskQTiwPppLWxbbk+g7lwzQsKzcNeLnZJx0KHcNaLUz67yJqWM6S2q6L
s6Txzkbe6QDr/tCYai5UX93gt+avqG7NFUSD6koEYNNpgPV5IXh3CDKh677Ebpx1nYW/Xp0Cr2gy
2fnstmVh3I7bR/5loGYWcNuIgdafV2Czw+6OpLWYUanuJbjnhRHvzHeldWJNPUTUecwO4br0MlXK
jbr/3Y96wVQI/FaoH4vGnJYG2brJp+y3M5m5/p/5PKAMpynkg8J3UEtJgCyWAnZQeUM+hWAQNS6Q
3S7tEVUwPIVxTjk7FinHUTBT+S+bJWuJhdPsWLPcd0bkrbstEo6COogpb14B6Muk2OA5bdnUpk4Q
zjcAChJfWwWw7i1EgAnZfQUOF5pg3FkFAkpetGASD3DDnf0jDk4xNtetn3UxcjXSveGb5jBGkpLh
pZEBTg7pHwJQGEmAmagsYTp/NZCHtevHCmX5BrFFPRQyVAdcCtJnDhDp55v1x7uKGBmeTdcoDKF8
SwTzQAQ56lLcbDaRQK7ezd7B04zrRo/ajuZnMSvSyYJTFFP9rLkd6t6fGnEw+EYPmFlu5RwohuMw
JCod55lEM/usayo1s7GNZu2YHWTKzs1q87pnXV/2xVwPa2XGY8GJGkdjW6VbF1HUYCsB8jNAUjpC
L0U2N0tYHh5q5pt2RDry+KhuoiwSR+K95UYjgyBybDSqYBLO763FaLO1X7s9LYwBDVe5HJbu2VQ9
wX8lqiFJE2UnnWC8dXBb9GAZNK2RTtVRXqYoKUWbxv6MFQh0uYQIclzJbpPAQemwVQGe1pT8IfOR
4i3iu9H/GErVqYSGZSInAuHIDxA2XawohCS2WjCUGrLVYo28oJg0iOXqlxVuojmwgtED+jLCRtom
Of4IyAOTQWQ3xVyws1Fn2z0HnQCeVkTjF21nvXSnIuxno8t3Erz0NPYujQlerzXnSh2kBIdSpZMD
kTKy7f2Ue25mMIhEDyhQ22DrFiB4OdugrcDbilJEKPlPHSydds+kCB+wzARHR0TjeoNP6G96yigf
84SV6Aw/QrLruFeH7+g1i7QKRoNxDOaF26Z74P3f6/5Gk9FYuZTCh1IVgQjQJGt5WBe+1qspyI/i
5hJaCryP6R6FniSXmXIUijLhtE+DQEFCgUSzUtmAM+Qr2lTVjGyQWGB5BkYYt3TXBRFdJf6jaTgw
Jp0AkzGF1G8ywIhCf/cqoc/H8avC+TbcCPEcg42MeFNFAvORIrKnxpTKM4XkhaVnkykGhVgg+iS5
m7gUdw/wbWa2XCKPMnQu7ljQhg4X8FsARjo9LWWBawpgifj1+V7GyxvE1HQfqNaLpvL5DMVUFiFJ
3WmG8Q44VnL0SLquFaMbktmCiOzQ12wDqKmUzOkqIAqBSv5phgzWekD/SNZ16KutHEgQ2ZuKSdsX
74lbrt+eCnxAJa676hD/KQ4Y3zZnc57Kx7Xga++eU9b6vTI6FBVAlpuXeg3JcFWRqWQQ/VU84x+1
QnEPDxlC/ItJy67J2++AT32BMlp7oNnKhruClwapOmOplK3wAPwQpWKrBzt6Iy4Nzjt1zh+oDscK
RAmzi8atw4cw4maf2v0WiQgSpnjWZ4s6rPY7/7aT/tS78x0w0np32pRvMNQwLmF2Hj7Mz0bk071V
Jifc9HoB8c9HgjRu0RHb3OD66do0RKlk+OysartYKK7YFbOPW53QgGF+yFJ8O1c9TyF3fgskePhp
Zx7GQYrDqGZHM4TUZXi5aUV6WhayWMIj1Ycb7Pg+d1L0WvG/b3Ts93kzFn7UlAJnXCebVIJ2EyLD
yoFAzQgUXSOZxRsubB2Eu/UtdfcqQBIbH8vgcF0ySYpaZxucTc5rG4AQ1fhpi6+XMFAsUKlOt7S0
edhq1q2M7ZDwTCFKjPZTwV1paSPYzvH1ypEJI03t6ZVlwWGaIr+QeOTgo1poReJJ2+9Dz85Kf2yr
IIn9uS9dNFcmiLddPrvd+4oLaOllzELa2VOyMU4n5HyqsC2yuyD6RoIUsBKTeJOFYHfAfop71l/i
AohcuXaMRgpBbfgRlVUVQEnorE775fHX7LcS3gkDa6wgY7jfOksESEGddPQgf+M8vaQiI41NhSJY
K5PlfIl68emZeoXgU2Z8OdSpLM3co8jCrAAauVL8TfjAYTevhLz4fhv2Lbsn6WwsIpy/BQWYGG3b
I/olC4Mp60HNE52wvXvxlKJvfy7JQPkvhHAF6N6HqzMRAFI4j6v15dxkgxmYGid5MZ/KtKtuEkCz
anYRpJb+k7CBZisi7FWYlHIeyyJsaNLGApJhHE0qoZ1sFKxGev9o1CI9tMFEkWvr6AW//UGExU4/
iRZI3guZqNNIik3Bv9VjnXIUEu26dDkUd/947ZMQjRfK11pv1KiG2VGYubR8GhZLgPcTryJf09mC
nVCxSGUBgn6+ygznvPWLB7LXKWqImuPZ8ZZRAUprql7Rttbygog9BcweTtyjlDp5c8vos3qZ3TYX
uETmQdbrk/LbeH6i41NAP8t4x6VPkjhyNE5xXi8/BQ3Z63Dq8VLA2r+FQbgQ2N57ydPX6lLmYFuT
ue6iLS5Q79rFf/aY7bI3DoJ+Ff+7PrBH6tgNlE8RlyJjiwkzpvm68OGKwq+V7VP8h+kDigWMCZul
tKnAr1Rf7ofTGcozgjmRGVmXsWR1xDZTDKhY7TrrQP+gt7Zg8IkBNEpiEr4AbGepAxYzhTNgvBsU
GX0iC1bSIhJw0jdApPVEvV0sQpoFlSSWz9pdLP+gQxeYftDpmApJI9mRo/EVGb1n/tUAmYWIvWej
nVLX4Cy0V3INAITCVOEk/tHIjWZEJT0QZZulPjWMUgaU0R7UKPhpHTut4qStHfleNKWs+/ZX94if
jUiSRsUiBae7xTnNVQeXXH7XRUwOZrD7N2he+jPRwnqRhE5xz83yO4CXseGoz7AVI0f6TmaW2Cja
LmfGe09ZXchikznSC28qiFEuxE5wWgy/b1Yl+F36xrMF6LqX8u5hkJsFJX/aLQyCnmEy8XnmiCX6
5xirOG+vqi1iqE5G9YVR8POxQAIPld8PwP/gswO/21K77jWcmotXJNr1tySaL/ulA8z9Ac469dWY
d5dhX5tEJpdzhqtkZgN5qKVUJsWOrHCvcHkQZG9q5za8V0tbURnTdW9n5VakGa3eBsuFMHgVWy8f
L7P3hDRtjmgRBeNjc9kpW8yM77fLbtN6d6UQ2Fq5RWJHdx87ikv+5eTlyJZA/fkNe5zuUMOHZWPo
ntsilScV7ZcmXFn659ErV6LIsSEEzrKPhAK65t5h9hpbNEPOENllV6qTAq02zJAL8Vt9rvsJkvtq
ZaYnopCHnx2L6kLc2AOICjT/7UNUyKgtF4ns50r/dmG+o6vv75vj7yA8ypJ8Z8aydARHYJw/I2mA
LckGWKM09AHjbD1zfPiWtdiAiAhqOfBaUSz6rwk7TRHm5FBP1jZZFZN6EflXpsVJPsmLjtU5lUWJ
Ihn93Qk/zmOGdFsW3rGnSHb7WnBc1v4T9WHIVNBm3LiyTVx/gXly2+BVc99mVF4DT8KsFIi+4YSA
pAf0Els6hGEP9d0IWBHYOIWd2ufWZkwB+nJPn+N55+01b0Md5uQmSKer/qrHOKkhT6N+uZMKpX+z
whq9CHSW/u2Y9WEbH7mFGoJhpjWsKtr0h9M/7DycFqnkRXxWbgvt7Cm5XoL67vzViO4jQgu65G5z
rqD9Nc87CWpV1WlfggZ4qg9NXMiTUBMwTdbxiz7aacj3DdhkUI55r36/rXcKbpkmYxITXtxN/cgg
WMbRGW8WnT+QRPs89Vnh2ujrC4Gbe6qfxjv/AC1yoNIyLT6Cy0Aqe61ruHOfEr/eB7smkby7Vh/g
r8+NtnewySuLQqzeEqMG5eVgmprVlcChcG4GjtgngixU6ega8w9yrOLo2+l001tWL5LZZn7hODOK
akyL+pcq32vkNKsWJGWVa0COhCzyanRBZUiV1pc2LiXhR8H25kOAO/4huM864kpv8SorqVAlcsj2
wk4IRMCfvPtIgitR0Arz+J8Qsxm1umJ4Sgps72zfpHx2ys3SVPwzsguPQHbM9yr5IuvkYizopc8b
x7Mkc+kKAKkZ63u2oISpbPk02ltrnGPzgVhZUJafxfqQBoDTDTKjimtoUpTsGUj+WJquIV2XSwqs
/FTxUIYrq1Arxip+i0Ia0+b1ouwRmVxgFOiCNqORy7khVoG7vBOyJNHqOkyykDvO+iYXt1Wuk75w
xCxPp50OdwTgLkncFmksGLMjqBOEk8sdBY27MZZCQqcVzhIz/LtPHrhJhqJCbhDnK81eYO0OTMS2
w48Rh2P8W3crOonqTpEZJeFRXbD3QH232e5hU08xUU6N4wnSSyVqMOAJ2Kp52xwLqr0Jo1xNSZzp
7VJgGcrZr+LWogAwLAP/RKq66q6mHaJ6DxRnBCzRpe7o424j98Sp4xfKYaUQ3lfyq4jLtf7IV9Xd
3YmVpSP8KHSHskoTZkaWuIOetZChmeqCpQtoFfZz7RkFM9homcsf2Ma/08yBuCtOBD49JqKHgw6Z
DafiXrzuFX3JXZBc62Apm9qkMCcxnGx4MDyQam2mi0X8Mq8fX00vDFip27PJ5yBkXwXScKU+vWi4
6EybRsS6S3k7/9k5zCS5lNA3DZOLwzE1BPGc4+935rn7CfYlnrNJWT+NomvOmL167Nc/eZj9G4Go
COn93OMByrDgE/mfeye0V2CTWg2qaVSd4/81NINGbaPFSUaL+nKxokeLbopel2gRHwIkDLjAebg5
WoNpm1wTUEvu/coHx+9SJ1F3bwxi5CLmIU96ZfD/Qz9u2GI0ElOaXDkFLYFuf+iVzbjhQv5wEmw8
z1DGC2xah7POsFet2fjDmSjDLTICSFmo6Xc0g09aoRWLpItM6WpCF95jbq36/6bm01+xtnFZEiZP
CRCtLQh3FE6mRyyZ6kommQz7TPAqt1Qiq472Y8YL0X2GNMsFiY+lQxokKacWUK6+fbcbRJdGzAni
jOnpGh7H//KQTiNv9+9VSgwKf0zfXrnD6m8uA6APsPtx2mj6dJzM69ChIr+kBXKnzQyb+baTumTI
ajKmubQv986vpKMPmz3gFpsOSR65wmsRiNoC/5IjMIn6KPSO4IDKcBlXpzwXOrzP8FtDX0hq+Y03
OsppE/906ur2L2ZLh8t4NAx21IAUDZtMw/ptunCAWy3NLjeSIRngJudh9d1T5aY2KvLzixv0H54k
hc3aLcladALB6T1aIdLtT3SU7cXGk2Gk+ZOBPl/fmm0JZ3xWbweMeDmQh1IjxaaNKqu63M5VwxEY
DJqNV7EupNltf8insyRAADhBncQjyZO+vpfaW24YBp4gB9Hnhs7tBQ9h5p+1F6mmGYFj1sKV/kPW
uB/craBELGPd5pp1GTzMDa8YXrByyiE1n0tDegK4D4j5I8gx5E2daKjpLonIr2GTzxkXup5m0SHL
WJQQAa5eoKPsUgZPjGOEf/mdBt7iDYNIIxFn+EqlpBj0xIBZn5V/NmsXM/HNRNuWzSQcjDmsuOW9
UCuqhpGvU4Q0/30aB3pcZ1ZjtdQGwYWOpCVd7J6HVx2mFhLs9b79Jo62i5NW3Zz8puQBmhG80H2t
VIKSxHuDV2A3AbL7vei0+nXcdl+3C6boIHUoSZZ9CvobNCdIOs+Jx9OyxNCqZdb8lMapUJRZh6q3
z/AwcwL5XyoWHFMICQFbgJfSHKapKcamTk4R32EOOZndT4Gr/A0vbvsyNXFnw9z5Y+mluwKxg13l
//BWSk1nYz1Jk9+3k2x6kfwKxD4L6OL/7tPvL1XAUN2rve5RkAWkvvjLF3FGVLILoOJa2BFI7taI
g+fdIzFg8/7gTleI+Hanw3ZTsNYbjSJ27kJVqj8cmj4mU0hyS8hsgQ74UWYpviEScUIBUdzvuBew
sCDbPldpVBkmDV7+sKxVoGBoeEZhBZfCOQdUUA600KjC4PBbS0O1vtQcSWsPXyE3nYhD8KZJmC+a
EckSWIRqzR7qkotCrmiM03I5hCb532OKp7Vpw2wH7DjYJrYOURaZ1vof8xZhro0/YUWQ0VNmhxsO
YW4a9fsvIgSwQ9fyKkgJvSg5VbY8Ib+snaFSfsXCDhQUV/HoZp4arQPcPReXQN4C3NE+nRWmpFiX
mcNrPL+/z/SP4uyD5grNx8m68fT/CdeKv4bAS7zk4N+R8xDweW7xd0xQ845to/c9JE/6KlD/KGB4
qTJDP48LTVErMDTB/z+T3cdcM7yS3hPeEQ7gqcZAc+fPEtIGA5eTPP63YMOUOnOA6d7Ta0HJ0DjC
Ee3IEkTxwNrq7ffgqsIvb5HQ5gXIYR9XGED3+HKnggZUdNYpmnRqP6D/6jgr9UwFpeaWCrtltndQ
N1KCYAnVJ7fVh5el/OqrKcTRWR3n2UUsWKCcOuLlzU83pDO/mYDMDc+AhbtOzf8/Sw94Cz4szI9n
I4WZWOql69j4XnoBrkcHvK/RY8DfpheuTiw/b/Toqiuj+SPYjUwX4XRCbEkI065CFUlB4jssAi4h
ut3qBQ8xSN1XNnNvpwQ36o1peUxi1XBNnHOvSwlTiM+/qvGMdS+Pl+JpzwWPf1DueTg7VJKFEJF8
dl4UAHfcICgGmitWQjUi3eoA6ZEnKJsw43KjPYzsQ9pxnpdrXi3ojD4BP41JwHbZEnun71xQPXoI
M11mVsc8D5eGJJkk8lrxP7OkcMpv+M/4gGEU12g2Ct8H/1MAkkzMeNRXN8kq+qimHZU5ynnV9o+l
CfE53Vn1SikUdwkx4JYfzE3H3+l4xb1e1tV5+PnR9/3Vv+9WzCmbhOkdxIlmoO+MHS/3pfTm9rKF
g+fhbsjTQo5QXhAp+576zK4LXzydcTtDFNy5sOyGyerQ3aWkE7RKOz2PzcGBCmLQtisnUO+VT5K7
I5f2Kdfvl437/oLWuoDQmMA46xIKUgRK59nC3ZHQBjdt9aadnR1nz+COgS2U4nygr6ZBuEr2wjPv
w72W00kCxmSa8B7kHGaSWLb/xyrRPQR6/NAg+pTYWH7Rgpq46An7THH0WOBdsfVu5XVTUYrgfGWZ
QpRJI5LF0VhHA+ZnqYw+gDePrOVgtmiV5B7zU4gEPnyJkqcJA41p7my06LIbTVsWSn5zclxjv1sX
BkenzxDRTszYtN/CIIu84t2pfSDaxWkLU7/tbw0ugiU3FiMAeT4KvuFNQpjdJVOoha6kiHyG5g9L
DmcPbzNUAehL7eK90pY46tiR3CZhw/GjhiEylIsAEj8mckAEYsry9Fuj2/PBEnabkajOcvbVuS0i
qSzABJ1rXPyPmyCDQDiwBwrR8Fz9p+WFd+Dyk3a8T85x4EzPH9EtaKMGNhO5vAYd4bZidqgnbcpR
qaPvocaBxgq5SSRP0HelNYS/6Iz4jY6ke2IBdSRn2YfkaKF/OXnN1dc/W/BYbc9ZHkBrxGLF5HKW
nEkZmxcaGb+r1yJlis/95RVeBhaIyYU2g+W4j2w/q7++BEuRkIgr0wdhwn32iy9bmnJEVIAE+L5s
AeYxHrHZJmgS1FeNHTHcE83o5rFwhfnBSz3qFBd+hBxVeRd76+zBDKfTI28P/PZIHxp2jaRvaOKZ
Q8ULI5He2DbBIGpKcvKwWxdBnF6cHYSxPrwzhsbj3cUEuonAQNyVp4AkzIvnxeTJGEhWlXkid/6F
ygkkuucX7U+Q6v7E/JVEaVQQO0/qPMkbTwQHPTRfCkLw80b8NxRIKZOByHTAhwaziZ7vFxeUuIKP
k6HLekVCB7QfpOyQl1GaV60xM0RpowJOzPabQfN4HrSpTE4ewS5sSsa2WvtFCUdh0aELidO85Gra
2YM8DFC/N218a6xzY/NMcPs5NpIFD5WZBYRgnurXDgTDli5blohLblQs21c5XO8uIvYJ8Sx9z0+v
LmpgT3z5l3nlJT6J0sdcVZbBAHSYgJe1wO2rBXdu04NAIv+RC80VZqY+li/cHpIAjt8o9GQOhEb6
Q/uq60Z9EA9HMLhFazLTVnkdE9PMYPcavtAm5pXPm+pGtSBCSKHLh4DYEsqA2sQxqlMWIX94MDzS
yKIi8KjN/ZLunfs1QJIaPsjXebA5egyM4H8TiYD52ayvXtBbQFNmcUPnjCDksv/u8o+uq1C2FMt4
nahfhmsjWiLyYCVIR3nKL9qbrme1UynUPIBpwRMRC4c7w8bymFxlRRxFLL3Hi6MiNVULBKmyvwpt
LtpefQ4ZeuKQUn5FGATs/AhyO/lU035qEbTKa3xCHCKhbbihKN1CsLHoeI8/FW6vSg2a2GpLE1CP
uY3mvLYNp2gC1HjkftLpmxhF/LdeVX4AhwF8md4LePKITdjMYCNLAZDjjNzwg1XhnnmTH0ODtZLi
sY/AD0crU0sJT41jZtzOIiOWzgqr/sYgMG8KHT0erGC88Iih6sZpadUkuq9mUI5qoi7RyLsC1ftA
nerFDOAIp6gdukn5zcZ4Yuu/x5tTAl1eGG7K/lOR8SZsi62k717Rn7kE4RlzlXKS8yOfRQE3q2Mi
5AtTzxC93nTHKE/eL8XU9w/gXfvSrMUCPcwxWTs9gdgL36s+UmE/NgYNlWjAor7TfpkPyErGdkpH
IFlDUoRw1KcjyBE2MyhXe49W38nW+bgxXx64YF6Q6bvy5CV+hHoBXc7eQUFmiFGq97hAfuOlHImM
9d5FE0jGYVs/yK1NLLhshJGWh0Zmc4DgtOrnOKsJAx0bT65cJkBbNKZEbp85mTfbHxwmav7TCfbY
//8oTxIemtwgpq3BqEYPF37O7pW+/bUL+3xBxOOmEEDnuGIS4I8GFA89CHzX2vo99GtjdEI6v8NZ
KjjVXeUEkZmcKLErHFeTbs7NS5JhhgpKXwMMNU5DS6LW8KzrzcsmD8GXo5RTUKzRwTpkr92oHbrq
Ylb1rpG12Dmw2WBPy7V1g6Ibwl+rHXguW4n5V8aIIGyXOxyeeHLH02rhmvD8asHQasEaHBi0G30E
uHz+/3Akpw96nvprXPoSQCTmpL9leDplxuTDdgllA4E7nDC1tu5OTpSXrAL1Y1LbTjqmyFUG7fTA
umt9Iby6eNgDxpGFrOJBm0jbiqh6p9lssthkCO3IGt9+DRo8AuYiouXzTm1olKGbOLC5VoIkI+Dc
vLiZ4Yhd1w5NZyGUFpUcD4hkquexUTw+lsSBdzTmav/lp0zdjuU+avxuYYJt9nSE1MnXerEbPOsE
J7guHjU9EGqIKZ263oaMQ/Gwy6I+Sx22uvh/kgzNvUuTz+Nb71XFpXvd66scwWy2uQbriGq1KRHy
vFxOEr72zQrRlxkxV1YzGAhXJ7ucDQsunxeb+1f4wyjDwyw5qJPDunV3SwLxBt82aznNkP4dVgTE
XnFmbKsG0SkeNus1VhME4WohYkb0a9KY/yKo1E3PfhZtRlAsrPuy8gFEL8goeAsv5maLA6wBqsX2
tK1sAB1+UqhR/IPThToNphpd2TIBgXIfM9Y3NoXJDG3V9hTosA3/C3837hgpEUd2wp/uZfZi1EcW
PRHNEyikAaKObMOKLU0RUtegbuAbJfVJZZtmSi1rErALUQAWPFWqmp8oKj97AM6bbAruZkn6gdjc
B0qESV7GJaOZM/QNeFTmtDRsy7F1tktw9YmyPPM3zqfRL8I56MelO1CwOE5p6mNpBQt8qDUQ2FHj
C4mDrftCLxTEtRFGM8ZsEtFaiv5LC4gFuj3zGcxFCyN7iZE4D4n5BwqTkthnPP3s4gc/arKe0d3L
SJWxbjLBnrmp+GejhPQayhQ0a4Ob1eD/7EcFGC5Xsm6LPazLo8/xq5CDJsvSZeIv+iELDUlspZcP
H/VVeMabC9b/u5vlt4uUe00vST1hAsXC3SZderiv1r3Ex1nOtzFvkAWd6S7l53OthuGNYoSGtn1i
FdcCIR33RCMblcSGsnUQQVvHF2MkVGbKZXhPRtaHUkcsG5GImtkjXrSxHIg8q8xN5JBEHFgw4n+y
egXAcL9XJ2CVYlfeut8RtqvlhyswOAlJ8WsrzeZXQ3WFNuA3po7Nssvbhh/eIAuGfR8HicC0bWUu
+AKAmkpF5fvU73OwWasrFRNo9OnpoLerE3rIdcX8ieRgfBfjvNO8EadOHSAL6hRHSI1Exs+hYbQJ
CARLHzsH6MGwN2axdfMEr2uk8FkoAAaLfN8UtKkknflPJhv57lm0huL4JSDDeCzMnbDQuY+82wLc
LyGNn974b0u6S81JgjS1tXcoiY/LYsJuZK5JzLelqiB/6+gS8ifPxUGm+0RPidBVxcvi1pTu/dBY
wmUAPa/2WLzFbECdg3Z1toEthFvpvHlC/IUJzmXo3g3Yhc+C7ZCm5muRp7jY7cubB/2/p3tw+bqD
6qQDjnOWKwR647f56ayU+m+cxCJXV2Z2fnRhB4Rpwo6imkN6tQNgVJ7wAEFS5SRD9LNP1yK/dfVb
60VoPfdwBrznqU5Nj+BTxNojyjqMR/SJvC+RUUemGRQE3jZRTw79PkQIolSQqosxh9Lx6jgz4OrS
bm+0vbT8sJjrqzZ/CPrOLJJqU4s2ssqiWsCT9RJbxBXGAxPAA/jga+3G/eHtVogCcHof0c6eID95
I4tnWo+M8Bpsx5NNNANflmpwfdpEXk7TgqpO3CTMxn6h1RMn8A+bQeAxTAcPDGoEu1+8pspeTY6i
gy2hiRipUDDnrLZJk6xlBv0G/APKAqNNB2kDyX2ecQrGMDWXO5tlk2HbMrCEym3Hkloivtbn6K3X
esyeCzkfzwR59ANfBaqrfGgaGkj0xU2LBIa2a+aPiqQ+Zzny//kFawEFruiZYyB0FP8JrjNQq6Qt
Cd5+yVYfbZyvcFhAzn+UyAc9PoIFRy243zq+6pozdVx9KxAJBAKrDnjViZ7qppWXfH4p0XBf/3xS
GycI4n1iEqeK/8Wzr1OHX0HNaYFrbA+CF26r8wCRcmCmuzO2r+TvZBHSchKjiAVnUtPl34N6/wWV
v4bmcVg9PSoJ8Sd6n1y1s8U60YYQmGMQHz7cvoq2nCIFzTak1Apqijxfb0cVvTlPS2ENyPw1IlSt
vrebhqBLSvQ4quFr47GxEQDlimtNeujsbRLI+ydhJsB/Bydk1qapaKDiK2VKG6WzZ0Ul/+JEakn2
N8AcfDiXdDWiRICkte19VU34lNbrh42xt8mWe2ZKHpHNP2ynhUh7MIlMtmQ+iO+XNE/o41kuTsEk
xTLWFXfsTUt6i5FVLOY4yxXxZb0qEgYpWAZozbZ0I6b8zgGGVdaQXXN1lwV+0uy8vrreDRR2HByo
8XyAqqEj7bVVAj23VOVX/0EJ/9y5/AjlpbGiBFq6xjviwmjTxNcx2e9wULucCQEF5YCyKWsa5xPp
9X65vlizHo11j2WzOJexhmgymxyPQcAacx+LcdYnTA9HHbQwWG/xL6xjkC8sfbEX6uotDJRS1dBg
S9NoEGhO/zMnI48/+ELms0iZPQZNQ4b7RW6o41V3MnVoFi6vlxSC9P+YUhfarelYHkyRfv18bbzO
OFmdwuwBwGlwKztmIDwQ/wMhuyL6vSFDUya4otZpSRSdG+A1rjp66iAMz4uA/F4G1cct5dymFk5p
BOBW2S7heSAD5Y3NZqIWOXIy013MleDMP/BiMg1LV1Xf6mzu2psFIvXLb/5tKKt2quhn2sjm1w+l
kVDnAxpzJiFVA3wRlLklyKNcTw3o5a1eAPUh9Vwx4kL9q2gCFCxRVjQ7/B+3avQcRvRcprAQEapa
th7KpkB+A5BeESRzDcj3Kghe3wx2MeWUVKKrSiQk95CTNTB242q/dqzbrIu8RMZW78P2yyKLrAtp
C+ioYDzUcSMYUrPtBRKimgmWWHm3wpBgTnYs2r60YCGih0V+b6EWlnJS48AkhYTrPbseE7z1phbZ
izCLlOVwftyoovM978uR1QqjvQV3LU0smoajODoyqJPYrf8oJKVeAiIM8PTX3hDVbU4nKq4A4IfM
QYks68r3dX7PG/H671MmQig5f1w2Hr3pzAsmCWw9pcTOLO7qX7navu95S1vhvkiKEAr+FfErgcFQ
uht5ZP5/uDuV+7ecVhUFDxwXfy4Fafx2F3I8vltCml3rx6bCt3c5pYmcrAVeMD6r8xltdJIn0qPZ
5uaaacqghlYdNDi0e1dn/z+Z4hsNZR8xm+DQ1G68SsvrmH4QYTdWeXsXtnZKdpebcQ5SADYeHbcA
jfh5RDdqx5n0+4Im/0dmtDt/8PsTCrV57UIul46DK11rQ+tOXV+d+kdKTUzgnY9kc7s7Fnt6ltTs
8gVicgwG4jPIlwwRin4u8U5ynamyvnwGLiHRGV8ZjjEBlLyKOO02B9NbM02Sa8snUa0v5HnCtcr7
sPZTJehyxbzbYMp2ziCfrj/6XdSUUeANKO+8vnNj633bvsYLuO2MP/Tu/gjEge1ptgWiJKdExkV8
BYMZFaw5Yl3TUA45r/9tB1IJxXlBSgxy38hhl5ZzVYXrnZ7yL/XT1AVRbHjxBH+/5y8OWQjMXhmH
5Dn/IZgdoW/nedkovEcncR8cVSBdHQTak+11XVvYOurqs86MoZCG4zqZxJWLbfuFwcmV6r4qxGl5
JT8XzFzXqezkKiFU39E2jbFAYCjr3H+DhClY+BhTwMmTe7DYAio2J45BNF1Z780l36s90f7ht9nU
oTQOQqpn49Wm7Vbn4RtbkkLATXrpFpLHw04pKSFM9dgTOrGEs4Ir6CEbhn2+Qmm4kV++aeHhUry+
o6Jg546+CV/pOQNkUxPQqE/78Fh8yHhAsGwIKcTPpQIjxb0Aca20F0PrbKTpiWeuwED4PDCz1Z2s
nTXq//nN5kZ7g51WwsZMhwF5jZAMs+tKm45fC6WZzLZG2o2c1iBBJdFCmzMZF2/ETiIMMYLYgQ0f
JMQgRTctVSfsqkUeRRAPv2MbVa23YrZmt6ksIGvPI3fRPUUndL6Mlqq2Sc0gnBIAnKHLAOqmsx2Q
00yaxL6nsOGmaScxa6TjsIkp332CMMP/NtiCNmebenpJob+OeFsNoxwXCSxNiSp2wN7YLTBLHpVl
nhJOP40tHSILm4lmpUkczVKw0WCbBgcmLxB1Ee+Gek95KfUqsAoum3o5etBdHX6+jXld+8rMGkdQ
z45vgCgX0x0I9GOtIwQoRoNBOTGG5dh2/+yKsuIHh3vGZ1OcqvNcI2V8FUKA4tBrkjQPIZNsDzgk
wQLgQjXAHBHiwM9a8OjpYrKb5p/YqpgEr9q+mdiXdhtPriz0mysEeHV9nOZ4APLlrlRpmex7KPU6
B8Xi7swJ1QdUts6HIGk6Cki6WC6qJK+qPtpWYdeo6NAWsmV0e/f4FFHHlkK7lQzGxZ5ZiTJ+Ek/s
/i+7s0QrHB5yQP43r/hgJ9SxMGEQVfH+C0Qk4XpSjTM0err1hdxA/TJMKtqpbmkZ7IJsXFYDdXh8
+Oia4SOJXJMuaVoSse2G2mo01we0ScFdnTbTrkEGzN5BWi+t+iZm76J/pyQIYO0AybPt8K1QwADA
sD272L+pNng1/8qpKazbV7TWw7UfTXsnI8vI4Qxlk/0FfvnGZTiEJkVgb0rCVOxWo7c2V2HSU1cq
bJsM3pfy3hX9eIGp+qbSis5vu3lQutIRHIhnrGJhkWZ+MaZnXyaldGAy7q6iAzc2o/v8yNoxYJNi
hJHu9JtbkSeJVG5WgDAMW2gacpCVzBXC5+ZkQw7xjXgxW67CdNisXI1Bp1yGN2T5171nKxZ6AFoH
RugBtmRuGOYC4H7yLHA38j3f54s4C7Usu/R1LovHVyN7pCSK6bt6xovD5t706Wh1oGuZEp0si3EY
Ol2Y11NVLOVr04wbCEeG5caZPdiiUs0/0kHS251ysUqVq8MiDDDFmSR5fh4q22Aq0CJF93iJ93Aj
plKxr5N8w/yR1IJ58pGeyl5c9pMkKHZn/QbIbZS1um4cjdE5TCDzjqkZFJGQVi+KChQe3+d4K8wr
XfzwSasFr71HQwwVZMd2zn1RXHKTY3D4xq6jZ5xeKq54I6eFJ0ksUc5gyySsQC1CaY3eaWFb8KeT
85XvN1y6GJa45h4BvTNT2Ef6SQK/3aFlkWDH69LDq/Iyd+8Gj+tJM74jLqsjn3bPLD0FMyt9Jp/9
Tov9vF6QQLnYx3iAjqtx2Xbs+m8GelPVQGH0gSxYv64D+l28Er28j1ElswLwV9bU63lBZwHAZNBn
uVjEKc1g2UAPDb0IkvVifBcY27kjFPm4ISPFVcEhQANNCiUYoSZCQbB5TWc3qp6yXopgoLBbyLTd
8tf3OXAW67g+NS+ZkBvK+4wUVfCdUrAJzhX5DYiZSbeS++aDgKaRxWfUl4hkbUOmt6F7pabKlxYQ
h/H1w5PzgtZh+N2koJsCWgNeYIlwultQhjqstmw8Ur1mLm4FNwQ2AH99Th8/YevjK7vOJk3FWWv5
vjiAat1/Dv4pEBjNe8qmnX8c5B3rpxdoh9RxtO05v48AnT0NfBd0fuUfmOfiGRL6xXc76ENDVFlv
7RVrtxD8pdMbHRLkQcPnbiKvuCdp7I3VNdx6xlCLFGfGAnuV0J5kXlQW0G6LadnuYXKJbeeU2VjX
YJYmpQVyrW9ZdP0UMjkcwgWeAYHXdGSLpppl38Jo6v1dHkTKXyYr18bhhcPoJbJLaWyczQtvWFwz
KEM4ItAN+xb39xYU2TudcyLXFCyo3Km0q9qMjV+cIj4R3isAqCqOucJwF9NPsXIizax27CX4ZDjX
rjA1Gpi/YE4Gc2WzxqLITu8614Z0s2SvY6/JIxQdxfcWCNSrjLfmn5K+66ATX8VGXg2LOUP/QG7h
bUaP1CWoCZm8Vhsr0ZAhceeDhTkosQbvCa6PYO8FDmMzH6GR08fvAOCFbbTZpa1kvuW6hBuTsFde
luBYcJ4WW7OCzsntxrRtEdIxbwRrA/X6/Od0+9FrvbhIV0EGLVaJAvWPiXquM+woisFI3sqqmS4H
ETMQ+Basf1ovBinf+fs7nDVB7yodBBIjJe+A6JvBPg+ofeVT14cRKrjzJPkd0088ju3Yl3LYCYf1
ybPLcH2XpLWgS85naU/8geXllDkgKUHA5tYQrow1R4/4O429STNGa16YFtuIScanWl/7YzzPsIX+
qRAdYzVUlBvGzG1pXXgnEeozxUwOlztKb0E4P3ZOn/J5vg3JPq293ltd9TwgROZ/DM6jT3ELheEF
s/AstaAXdtUc2B3KfuY6jht9i+BRNCgbV80hmotHMwFgs9ASJuq2Xq+bPIobASbZA+kRGmzSVZS3
hkFoB+twX6bLP/qjryWYHkPKVoLVtMGFcfSF09/4052hb/rK7jbwRqEOgYKoOGKOxqM4p76TZRza
FoCoBGOHzI8YLSsoygVbMg1dxXu5m4WuOsfEyncoiaj9+F/KnPGs9K984u+uSNKuWPzcPJWcTz65
B88oZVbXyzCt4sHpYoxdcR5JQNx32XFKF0Yf5MVKco47Plx5p8a1HJYcx8TqChWUddHbqfT9kBnc
1Rql7vB4O31rtDAQDVBLJE4jku58HvRHRSx0RN7IGedwICAZ/JYgpNForKd+XdLwbPxxwI3369U/
T1UQZ1KHyCt2B31hTEaZt3vahPSNZv1uwqu7hs7NHgBhVvT6QnM8WjKdDplOGdlOo2nE/PFZZxvH
sWQ320gfm7++F8fMrJ3D6E8HAMoSIcqI5a3HM4/ZqXmbHcRZpfXEpUV2JcHTzPRe/lx9qNChXq/j
qjuQsqkJgMy8aa6P2qToWBN0NRpmO3cRpeOcHkiBzrIB/odGoCPkCXnIK0UMWSA/SvJxS/j5gsXm
hx8FpRwkn0UjixXn2sjEKhnZplrZIMjv8vY5kmMT2T4FWwdaIyUezylt4SazD4/iltEJGws/vTdW
f7zwVsD4WvJ3lTQfti/ojU8SsxkpZytBjqPtMAy9pPJ2d+xfdpmR/jNo8CU+krSqVPVAvswwv1VH
HAZ9LWPAMiEVm+qEC1cbdrT5o6sTN8dQivi3mMQR8m/78CaCN37h+Dnodnqu/n636LimMl57gybt
8tjY95pUR0aiO4KBzgTJJT7v5GkfyEqFcx8lzeyZ7eY1WbHEc48Et+fqGW9c4l+FDIm2Lj0Tl8yI
mc8GSVG7fmda2xAYlIDyBtnDlrOgD5kknu46SU5qqKA2P35niH4fSzfSHq7GjzE0ZLy3oj4qx52f
r2EM159/j94c8Xcc3jHq2MSoPWcdLDpXuKmmVqmgT6YBTgVWoFGpex7ABi6+KXbT0yUIsp2pbJpa
+1tVawSVXjKHUsYXdBugdZmX1YO+axPt3XuHJ7tKjje4rNE4x5/GdQgJGOfZ5H53LA5yOUGHWFAA
OH36jsasodRhouI9VaYe38kY3eRqOaLLlmmTfGXaCOJ+5OcDD46yCASGbQwLIQB3Ga2H4Tr/Tft6
1feM8CwT+7ughgSsAr5NQhwROw9Ast6NKbO70zAq83gMR4ZzOB8xjAWLjJRaNXrT/Fyy7UPUiB9L
9rx8lPw+Cu58W22Cu/9QkeEBIn7PGlZ6aAzTnO7r4U9rodOPXKBp0QHGC9bsLZ238I4nYvDAgSDv
5ft2xdVN9JN8aOBsyqFl5iEYYgrEVDbzq4E8eQLnLBl5lmmH/THSKDvZ0TPltEZjsnEd1Y8hCazP
xb80jdv7mWe+7c7R6z8Ey7LL65qEZd7yUBKkfyMLGPLn5kl2U2oebAEdX7oraJf77bqsDS8u2OTh
ND3kalt6z3LPWMdwtsgDuOYZYej9v2BPMAcP7eZhQQvf4Qc6C3IFqQ5orTtp1x2HwtKQLSFjZj+8
Q1aEbbM9qs15T3Ckm+dXNh6avl3XepQKwqd8Kpz7ccUalQyGapZTuCOXaCU0QGcKq3gOMOV3g3Ja
N6Vau4mroR9Wt05+Tz2FUZCbq9XKQ5E2jKD431baKDFNeJiw6jLdIq66kdv6swqAFqCPfH9L/8pQ
aCRW/hi7w+KNsontCXjjCCyFun5KZTUvHYPRfdOJhbILLQfXss4j+d84tKjx6gDuvxg0h5JgPrC4
2WRwZ7v8gbPB1auOdbfq0x+ZyFLZcVlHlLy1cBw/O9Hl5JLlc73+XmVRgCnoK48FTi2A8Z6yFfTT
EQEJbaIumjU5KFlbIJBgdUndLT3OVppFHIjwJIOHz3OWq4smY94Suks/Jx9U0mDxbxHCakFmrPj+
OKOGOEbvOLMm49fbRpEHv9vxXiR/IOGDrlzd3aDnlQvErHjNVLcqwWqqVzoaTK3mx7ooe5ZNdgEr
f/iaMP7HpTaqvMLvttZjxZPQnAcbL8KszGVY7khex+ya2xCyMNf3galLLYKRKnKN1Xu56fzD3Zy7
liuQtRu+N3O9F+2eltSwvyNB18+yCTbHNNrKvOJXzMmr+1uswwMoxMB4NToGncqrgGtX9Zn6y5tL
DkvMOpJ5P9WsXY80x4abnBeYACKUt2MH/IqHXFHg8vfNanH+MRW9KAao6gRPXiRpM5CvcRyb7H6j
p2fpYJLVh+zzbX5RM+foE28BTtC030c9rHBlBPD3EB0Nj1ya3ODiRiHoNyZ92Hh+rsWl8C3KuDti
slaMBUNZvJI5uXcpohZSsiDRfn7DbB2C3S3KKOGlRYKhGU0q7AUOgKeP1FPoNgKPvl7fW2SbMxT7
1P4cGa320xx7TPixjaJvCCMnJJw+uQoGtnYyZDWf/lTqhXVW1oCx6gTcSxD+i5pnY2Foyq/xG3Zl
Rw4zEJN+/LHXvY+r35z64dCcwS4dJiu6IstzzTMnf7p0TIvgaosLvgE2+iezVAkI0V3wG3+V31AT
oqpPWAweTdZCL1gQgqrGEOo/JiFBWK/JEjvAGCcV3zeSE6zr211HzHE3V5stAxxFXVJqvWNtXCLk
estnZkivGBy/T6po5DcX9Sf017RYV9+juy0+S3/iF2yXZAMLOgccpmsEi2Q+wypk969lJKR9SKza
zLxJ07x/O0Nt+HyOrW1DD/XBlpjrEhBZJmV8F3gY9i4Drr/Bhsnskvun5RLtB7qsMWkk9YcmRpVX
BliUCnEHZEfddEUcTfLwl2Gm2KJBak37TFYZIiXIfvDIITExn7QcQ3l2gpYW6BnoSWaKNXKjB1zP
62R0i9FkutaCyjNz4s9q3LeTU28SuUcuqgHJ+wB8oIQ+7/njF4hlQdEeBxdT8wwy6bYJaz+ec+uV
KDfIKb55QHFqDJgn6Z6FeIY6M/SIYBHXS5EiG4WJCubMXnVTVTGEZnJucolGAN/7v8Q5Mpwkp3JU
Ho1iPAu/WzewdWN5Af1oFFnhiPCjDG1nqOhWRAaleyWtH9Sd8LBFwGKi2Jdmk2LvtgSrBRHXibtK
eD8qCtlGrUX6UdU/ig6Is4hSarlNUHXeNAWqdLPzqXMahYTDIzk1hTNFoAbDSxQBh6siQ81Qzh0d
pf8FgsDxFURdD/yPia/pNrsoxzYOkhU68gU6GVGyoG2CwQBRr4eWcT5g+RkF2fHm40/VfHv3kn24
TQdC4Jk0WYT3FZtzRthv1WeGfAOHqP/hZZFSPCIGpMTRl2SqPQ2oXCN3wqjOZlsiv3IPXXvYezaw
rwolPknjqHf6Q/W5Qs7Lr9mLaZHYu015waG9mHCuM0E1YGuZyOujGtjHQ6dyttfGO+UIq+/BY2WF
6EVmqUgrkrIZOCMoEqkQSDewNvwDn+RgWFDSMKAXPj7mOt9R+W4teRs5o43vNpoxOyXiZiKbNods
BSqnnj2kxHJx0q17atbN1wmFvP6eSbPcItLDZFK0OvJ6Evfaq5uOd4Yx3Q7krqLjm67ITteh0cmy
QktCAzkrQosNohKvK8ZE14h064ZiuQ6U7LiSf/n1i2ta/uXJvPsQWiZ5ZiwDERKTsKfRa0zjruUl
CtL4xUJniPKuZ7coHs8CvLc1AFxhkkEyCiKsv0z3tDvvuYuq0VAIYRizTudhEtbABx2opwb91b5x
DIdM6AfUWE/Mm/Hb6SmLyqgig4kfrFmOSLkGq5m/weM7Ww9GsyNdSCIHBjF7FPzaeTATT3xnKXpq
gDL0GfmDbu0RB/IPZbxnqRJRhs4P9ekZyNzDRMmoWPUn1F0f7+ykwQTr1KcIfFulrnSY52BKqfgL
8K8O55aVLn+SDgvdtnhYUer8yi0dXUE2Jw0cH8zbv+G6y1lH85IcLCJcpuKdcIoTR4OB8e2yCGiv
MpfULoCRtZQsHOTxF8TeF/YO1DpuM/F01M5vbh0GlHXyLzexpu+4KLAlsEcoTzvsVndHg9th4bPH
/D2vQYaSu8IL8a4aciB48E3EESAT+/oPXkQGxMyJDlucFFqgBI0r2W8luDSxLRu9JGo3Fy0wXUts
5EQBxME1AmJPnY6WRRwJWB/R75fPjCNYPYM6QCxTYGUTGQINYkqb8LiFWUVf70qR7QzulR2NTP5L
bduMAhgviaxqtB0zDIE3ucE3Wpbq837hbcnN+c7nGuoKOzB52AuPofnRNlo1cAfOZ/rADVitiVLC
tqCErBKjBMuVgICWOAAYf/rXeFdTF1q99ts6LH4zOJD/mLgbaJ/wOjyu0ZT1YB1p29RUyxqIbGL5
Op6IZHTx8/Bni4l0P2jBb+1xQ+K91uNTj2czWYZG4ry6ipnyNZaL4/hy2blRtb8XEgb1sSPPy3Re
SBgYWvGfsBd6CXRJzT6nF1bkfvxEF7VGnYrIBQn2PB7vB/iBqoNMFnmzHWGeS/zJ8wSW1tveE/Ys
pObQQL3rYGNZNYf55R8+730zDekBsTMOsEckQQocwSTzg3DZFDHdAbinbpiyoeBP5uN+wcJvDDx5
ebUEXlTWjboPJCuCXnMUzYN2mlq2PrxKm2yAhtXb1P4unpy0wTcag46Evgzsjuu0z2C88GPd2fe6
tGMYzivKp1yPxDNokq4tRIhAT+gRhhMmcbyDUtA9QmJI4fG3fpiZWToJ99t2s45wRhmr4hbrgodZ
VNOuUIoF8mm8vUq6nfzNk97rWiX3PDCmUOu7GTY/hkmfaSF0Lt2GaDBOwhNGBYFIzZakG41svrD6
vRN/hxex4b7soZaH8L3Qh93oCFQ11u5m+X4Mif9jhIkwmwney3IqFzUAZC9LmlKRMKxJmky4HAAf
B8r7vs0oz7HWsXPxAan9KTCAvjK/7zP41tuo0HCU8uJtHeo+v7jHJNazxmAS0kCv1UO0pYYfgNjV
PsgWWp3VK15aiUi5nmM6S58+ZPL6cDcMXqEytomZtvxoc1HtGSZGBSnxAu8Vh+DCek/xjs6R7+Am
h2JKYMJWMed5r9lY9BlS+ZBaIYtifHe6tM7rPsi9pf9miPe6XrxSQuMuEQtXb/hhBDLgYdGjSAQ7
0kyzSiOEKTLRW4kiGdFK20cWwsIEluasIE3mPXt+HJPbq708WZdrUuu2bg4pfVzZQe3thYc2Ti3f
IgFCPlFlJSc9VvNM0b6LnkqnJnpSjbNe3jdTxEifxA4urf4hZ85wlUpxgc2t5EfOlhsYXdhH7evL
4gI7HDNUqx6rHZnRQz6bEwuDjKahC9rd/yMEC8jF4WYV8VRufK/wbjVMJd//CsCZhwCTFb9w63WQ
LRRkcKzzL17F80dRr9N+Zve6MaHVlN7trZTUQ1tfA2kzccwwAIWNSlldR1OA8UDxn73jlCQZXBJF
jH0eyuNfO7FYDpIJ/88W0uaBB2vJTBhF6bJxfCAabTS1npGEDEww3btZzKTY1jl+fNXS5REa1cYt
iPH+wss+fH46QqG86JCHQMbw4Lg/i9XKQosn6ikruVTc1e6MuDcE+zyJ7z1mS3Tt8d6PYN3xI/dB
7mCtUaZ0UuGVKpD9skGAFPuZZg2F2/vxoxlYINyBrFF4OrG/G3Gy8NZNHlFc8nJ/FJxoXYvhIpDl
UmLS8lFqMoff0YOqavkaycQ91jYEuUE90q7YGdR+8Z8adfdwCtM6kkqxPe8YqKjadn82OTxJ/7ND
JJdl4kabzUg0xi+k6SAATh+oi/LqQrLHrZchZDDEAiMGx0R8f/qiISfg2KfqCh+U4SWMfqIfrG+I
Td+Fra3RLzCmRsZ4EzrUEe4rJ4UTAYFjVg2ODgnFHlOGQIhNnstBUdT/Oe1cv6eD726uqrpHL3f9
u2qDygBGRXOMHh/BSNcqHfHjXgTZ3GuJy2THjMOySWj7nkw1FupSNB95v9aX9MkeW2QRGbvuDvTR
bqUP8AqrWn9c/F2VAsNlcSNb5iEUizTWiU+5iqBgwuW6h+NtHzLlRWvdo11Qdi0DQDhkGL5q187y
tmh1paMZTJ7ML2kET+U1ZTcoSQ9jlLy7gD5TWdDHoOQzFGASobCPVkYUwzSU0QH1Qn8zlaxawlCQ
rvW7K8z1jZR/juV2IR7OzHpe9n/xBMXBuyH+5MdBQC4vMWu3IjWlwOUfVOAEukRyniNk1osrg2Hf
aNMDJkheCqzPKABBiH+uSXbdYNJAvnWL4/pOsPTrTxAyDMI0U9k08A82XFZVT12p4xH2dByKxY4t
Rt9hv/9NYQvxrU1YuouBXNl7qOVV54urAOs14aQj13YzaUTWw+i2P+myJ/spf38cZMFlVwvptD0k
wx9FVeOOaL8m96IqnrjbZVsiElcEYxmX12tLQyzHLdiXNk07X9zVGbYt5LYwiu6HmW63Ypvicj0M
wx6reM7mOmQ4vvtrVxaqdzK1Gg6SMaG0XaWghQYMfb03niNcguCJf8aQc6Rcalw54W3Y2fI7TP+W
31nXm5B95buaUJNpT4HIAeifXzWp1jICfjkKfPCmDt0LrIcy1qA0P4WQ3dontJQL7AQUHWp5M5ft
ilNhJCaiXOPGLokfvl4EMiApiWVaJOycYMyV8o0B2i84ImZ7R176CkmACwmlbMGWGpN1OkhDv6Cd
gsmeP1RKjhqqA/Vf1wKmXno6gr0yUQL4l7rd/Neel8GTbKSyZesR+yK6ztSDzzaoVLwaqbpFCujv
eZFguy8S1c8JgRBFZh7e4N+eW0g5+DzPL7hSV4BJ1ESyobPmdldiWxPYz/8H+Xw7mL4qnettVotB
OdKy3MEeYkaiWRhY1eGEH0bkqxqb0r/4IyklzhdDkx0LlZ26PYa+pZUpcHGtF9ypC0V0AamTXJF8
lALEzQ1+OaEl3bPiLtDgQ0kPWJhvEkMWg+c77GMOBgYOCmSzg2UImXuAU7b5GMpk5yMHs7RAiC4f
ZflrmEDeRkNoiynr+lZ6X3jgKkdZwgwuuKpfMcxeKwJbHWHFjAetvqAU5p//QagN2vrNgXC93Sac
8NSekh2omndWATy2+7DvPmRsO9lyJxVBa6T6rm9z6gjACqDH+m/v6cvMAlMaiV48QfdLV9x7Pjgd
pxl434vj23YuzHWS4+JwK7aPB1M6ghw8HqZPOcwI0hj5XJRvmttr+lKedB3dK18PBg8tF97fCw2v
sUQX/jOROyhli3X1V9hojvSATevEWq/2GKMkDtziyeWQ+EjY4AZm/EY0CPP4bK+asT222xt8ffE8
PADmPQx3HdJrKLUe0JHvX3INcwEUuer0tx2IYemOTMfsWifuAdYgQaD+M3+hF/tyes1Gl0gybwyP
d2vKCGn4SHG/iXe4h3ePxjp9ABHSCg35SM9YJ321tPUTiG4siCkv9jaDFZAXooKe2oxmu8DwTyCY
Pph6YNfazAAkVqKeHP9ouQUJFsBDKpfBOTe+/A/HHjoTzehuipTGmmMRmBZkH+4F/vsSPDtUzni2
4E67TYN3KRXMtiEiv5QgzlXlJVzw/1rwyX+Pc79ysXHMQXhu7BISp5VSHx4jk/0q8d5/TL2DsgTH
f6nBxzfi2lkOcotNnLUQ6ZnSsFacPa6o9jdxeZ50y5LtddvS1Qxf3gv3jybUfRV3knRHkwzKIV5E
6mDI57j0vYune6/xuG69Z3Hrhyl97TS5AIVs7SEKx8ELAO13t3qtGjqWz5iQZc6hnAgY8sbyANs/
x2z0rZQCrndHmshayH+FY7U36j35PCdoVvwclyp1MFNtq6Jah3zM6n+/GdiCOlW1NXLgsTZQiKDV
pDNrJTGzpIHGpUhqu6diOLqQ0DgBi4e0iR/L8bGp7kudflmZtDPaI5JE/8ejeutk6l+0fpMgGudk
9ssnG4jWRj73BbsLtvG+AWzp5sUk6xpSrHP3DrEAo024qR4EuTarVEbzWdSvg3C0LjlU34lZMwOn
aAYer6Diav7AWalVbWOZclTr0g4Yl8uKfi5yEIVaOB2YrMs8graZzbmpzBBEpt0VnDqzNuBVUbrc
TkiqHM/Nji+F+S5ou99oDkgFGZfr3HRWukYenSqUEUgDWcjb7HtORKY6PBlmhL1Bu/phGiEzGCDk
cRLXryaOw+//PHodQ0kCErKGHu+sFYSxgrp+EeGKFt7FNL8anGJ7jW5TkuA+o8h5k26xtk+sVr/l
4+OqtAI2jdz1hKv+VLvrb4PGJB2Wnm4/OjJdUWnaOAZ8atxbC3ZOc60eVvWJXS4idu3tGjoVjRHQ
KSz84ZDtgG5NxCWb6U+qYDHv5HY8K0d+JjaLXUCco3nS2typTrxoMtwyAwTE62L8B13TLqBApyga
WkSuj+c3UxrqJQ4bpgdv9KPqN5hK7ThK8SyLktBGIOjIvelG3vE6wDDUYJuIRekCMCfhvyiSOlBe
FDIa0U/Nks0j/dkADdFqblJWHBJ1qpBpMMJeQwlvoarIWcKgmsk/x2mTba+Ohy6SiRI9v0bLISW4
gG5fy7IhL6BwAACCPDMsWPSqPjz0UFIfgG5yYs11eHXdQArDEv7JTU+3nO0yp+C0m+44Dt7/AUZ/
Qma0kpEHL0sRfjb3uBIA9sxd0nSQN2o+wEU/9phmgTvP7WW9q7v7Vy7YuV9SYbpXgp4cV5fcTcz+
1ohIqFaB5hDL/CeBul+jn7U+aAPG+EJNraWiZ1y8jkxYUMAqT9Zd469IcBF9VU3tbirxRiOaNCXP
z8Xx9Tx+DYzP902Bo0xTYVi/iukLfPZv/B9aXDmlqSh0OywO/WDL6nevtyscgHW4YA19hOgpK7KE
fZxDzXGBYiUA/F7tZeUEozzgQe44e58imx88egZyaHO6E+jqm29tJlU1vY8K0TXEZppngPctV9Hh
dpmI8fsSdB/Wb7Zo3TUemveQFkTiFH9z4dnGl6jrw6Ge8oNjm++j75HwKCGS4FCdy4bhKqwcFMn3
TD8OGMmbun0iaaqBCdLo1F/SjGXOI5i+pyVGQJKLQsulkbjmn0/0DINw1EgC0xZ/aJkr038F1ynG
xGTuQC6vP3lBLO00P+aGqFMvWurSwnMlomqD0m2FtrcE0uZnqOEo+LvHjMKQ6sgpTjP25wqENsYB
y/3GgURj3gAz5p9GHRuGOxLDr2u4gleZ5pEJQTEVAhXqDBsw4rquueqChXZBmNfVwClPainDSBDH
VI/zM6O5yO64nIPspHqljLOvIn08akBtquvzdiHbLpUVbSekfS58RTieDwrLdQnGgb4pbKUWuqvg
9AbBnw+EN674NSdmJBqKi65EyUq2Znu5ghOLwYRTQUKYgMaNlEhKLGmyl18jLB7PMEbvvrGnYE77
hzok6MCtkL2bklWHbJDX5ITjq3h64kAR0Wj6+jo28utFeF0HmzRzUtFnbYlJslk53KodqR+MZ472
NFWiSrCuzr1nkpKPkLFm2hU5Z26y+Q3nfnB5MkyR91JnFnIdueQEWppe0BdPI4e0X0aPtGBUxM9p
xiEcRjWZ86melIwkAHh2hIedYOdX//fUuzlDAAp+AV9EdYdPZmUk/JLHLH18nj8MJepuoZ2P5ADs
rAdZ8HkUxrxED0cKkvOc8nCZ2Hxx9AFcdGQXU683/CX67qnJxPO0C157xxIkYgpMZWg4wFs1t6YO
ioUF021GMwVcAp/Nkd2pHTfrYJpqm42xox7ggPR3QTZBywuaB0mocKntdn7bJZfr8YAnuwm17M2M
eXNZcVqsmAjRr37+0ZOF+Iq5EmASSnJFE/dzWy/d0n9Ek3zycWT2y+8YAg2BMtmBCB+Nag92G6O0
soDeBOwwctUHZOBtSK2xYwltRmMTz4HiZ3a4pWTgyD4sW9q221XtBQ/jzpmjxutaySBpX7GWPMbW
fFzFx/YPe6rEGSVfq0xIQdHzEOVWvIT1udRsnAbQh5gL8VF2tg66m2Jj+gBwtOQULT+OH6RKEZQS
Jmn0rJEZFKSJMXP2AfyTSbrhYXdwKvQ/2WDEU0vD07XzKfq/2atXOaToKS/H5TJ3ZWrAq6ulK7Fa
sluUmjvt8DwvbkeP/m1rBONpEp0nFXzf8UupR98edPRU4x0YUzXAkgJzW579RxQRKJit3de4BxTi
NjXZbxnNeq/1rjpjjl2Xe3bbW5WNFsNPNG8czrPDc0nXZz4wGrDjaGNEEY1fUrk9WRsuXqh3iTDV
WgQnU8E671kmlJxBwCzLKQaR01ppBCeg3FHW0NwMUx9OhifZgUgT7T7IKc69+Amn1P4nBR6EjMpv
mMmqE30sX5lwNkolN7Tyfd04r4yzMWmHW0SEBfdT/yDkLH5twjAyF6jrlRyu7/5+ky+rxDDh5y3y
awYS9cSMYKb6GTla2Smd82NBOlKtNbRLT9av7VJPIGiO6gO7zj0YrnWiyR5C7qdBkVow/tI+t13y
x6rKk06qEMFWV+6pC7i9G3pWLykDYFILSqAtFcOXWMoyuUmxnWi+2alX421D/7xHN6U0No5TQRd1
EdoXSrFywFfoJQN/q3EZL/Lfdp7qybqreXj/HfJcTCLyPx/5p+ckr+OTiJbu2dGVBmvVxUccAJ7+
zxQ2Z2nTd3afCpV6yDl6yAECTJ+ZyF1Z7vQlciAEkgDFa3Kqx9aZjVBtRNYjXULfKtjV8Ggu1tbT
w4W7qjX+MG5oiqSj48I4GPu5qaJ0/JMOv7EuEw1vFb4pYaNeZVGxSz9xUA6JRDHNGGYbtERk3XZq
tArO5Ivi1t/VTA6AUBQvZHxLfgizlkZuuexC35rZVnhhTqj33Dwaex4nBCk/mUVRFXesuY3PXt5m
OsAKKB91Fkip0KRW6SV2abrU/i6X46IMINlG5jjXgTqesmzSIDX5r2sTtzdaNUy+N5L2U2Z0SLde
DyKVIdUDEwUqW5Z2t+0SlDe2pwpoFlD7+y2GSXchrAfVjEY7WjUKHL5+T4B3GdQch0uQlu0sYwoQ
Q9D89qOeB7chWJWMzIpO+4bU3xJUNr0MHhCf3L/GtC1DHDvLVhoAuD0c9iWfsnjU9AmFhs3uNJfq
sTQKmVTbZdT6mxiNEh5HrilXCfswg4GWmWMo6k9f4WwDkf6Qr9eEUa/B5vY10AyOognDWPVvK+Sa
RzXL1z+1mY31ZZWbV+t9oBzCLCy/FqYqzWDog5jDplOxx8m61w+z0v6//Ve8VHwY8pmYybt32EDG
xgYronYkyg95+9+Cok1XCbzLP+3wA/Cg+pOmMGEfq2qf+zyPNQ0mkC2wkp0gIYEGsEUkNv7v+LLj
BY7sCOM+6Q3s7TzQ6qGxlVJqdOu7smYTAFJ9b0ahPCo69RPTM39dSylVTG/WS/tpR8dVxN0C6vtS
nIssxQ3Y/zo+5gtAulraVLUkKDh+ppqhpl9XUgdWbBwde1bkshe4dDu7kdmnzwMs/9bDHdErCU5V
hG8p1pZ3i4rDyz2Cze9Lig4tcKpFxzjs92EXpnylNKUSdS36lMDyJVWuXIq31C2xY4aB0aTqH4l3
kaVmcb2a/sqOLLENk+DL4wc2l6oxkUyLj/ywFWn8ht3Mr1cmqB60Ks7Ar6CWcTeo9Yw35vbmjkBt
fKXFqJmH3zDG0kjmy4I3BYd9yLvIwDu3Sc+9eouE3VvroxVP4juwpCs2J1fWVz6kPkiPRaQ4BGB7
AVpO8ywrHs+LiuTKphEISZOkHi1onnjbdvImPgafhB0yWBh+r+5rSEuhmKvdAHPzFj/c10tXyFhs
p4hvnKGa4MLBhJWdnb+Bjvt7NXx6ZSURjiZUv+5JCuWwUUjBTxj79fZIGz8x5pSIH0saeL0HleF+
YsMWvID5HNswWmamMGHG1+PnjvXkpJgLRoLMVE+SgNCc6kipLW42DEzZhT4oimrVeCGSR8iz9qw3
ba5y52VAzAt66oc9kMlNCcawE7qamTj92NlVez83KYpIYSWgOtCu7X+sZ55NwnDO48oUzY5Rv1BN
7z/stnRxplSHSlQuyeZ5hQ9gHby285ylQJwf16EZ9GOGb6reANDZMd0UVHpo0+UOR0kNLRJp3EcT
jleO2bEfeduZsbdabo0QfYpEUW2CBfmyS+f/Ve1J6vBjALRNA151VpUCbg5fcIC8BUqjY3usZ+45
vtMDO08qMt1LSQqtWTT9dH6p5r7MR+qJSy0T/zAf4fGQCj9MhibMoHVUTY/Whcn4/Il38RfPjIcc
Ld2srj4eJpoFpzPaI8ZI8Pv7yCB3ESgZD8KdNzjzlCv5XZeHkraTH6asKHtmb6qiLEZm0bHEZrtf
JhLtRrCiWjVrWsGYoyB/6otV/AvEfFuMkwWL0r/LIRUB1eN1GXUrx6keSsFfzaXJtd+IZ8/3xw9e
5dp2Dd3ZKX0njriYv+V1EDi4zTCiaTokJBcYlO8rheA/HxQTEtDhVPVUBVLZfucA8bG/QBXJOUaM
eS+VTN+VeDyutKyNmfqEpLP4l5f4LFJg10qEDc6llCYu+rl7qZb6ZgZK8O5MU1NyVacodAN9eAzX
vMNKD4Y8Sotiimpy4NFFpiwl0gjPtrDoU21wTznLTUckmcaToumJfM2O2NnU/gQA9l8ZE1vkeVs5
nk7T02+PsH7eL1lmg7oCMefpkhKtiYvCn0xhucVrnJCGC3jybaSm/TYjYbFDED1FTY5AdukY5eeu
UTdjUzmZlNSzoSj/LLC9nT3ZUvGociKmA+rf1gS5wreG1S8eu08wfKuHD8J7lUeDXo2WSO0MbJgl
ZK+gQXzksiaVP3wyUnpjerXLQwVhgSkP/9vPUJQsWBwO4lpfd2DJWMK/c1OV79iBaVftimEjE4G0
/04W7z9T2EIj9mFKx/gh6e1mn81ML35PhPH0a+aymK04yHU7uNfGSIwMONhf8jndQn3uEVrf4TPj
BEvvxgjOUiGsL0eSQcskwZPzYSo4IO9w2tH20AY0QFnF9qTOwGz4K4Qs8/SDOA/U8VZ8iftwqdTO
H4dMJRhveVMdDXR5pGNQOp6UYdGsGTf4ydBLKDJU2sCqow8b2SZe8dRvoLCjyd0TXrSglQeB/9mi
CjTBHvz3UeYOlOSp60dZ9Mcg6u63J1ZI+3Zvl2GmZ21/n7OfJ8+MS+7LJTmGcoA7WoD05NHpDJpa
6jPvY3Ev1fcZdLSy1EisgNxuRHTSUqnvpj27E11JntIlpl/EgbdoMhvl4Uhsc/ugfFv4Hb0CdWW5
bgADQqBp8hyMSsQCccJpi8bWpnE4vvGnHLFtUp8SJwnqWF89Tny/cIU9uLciXvogiYEvrxp5zi/C
YDCf0o03M/y96+9n47zu6qzQz2ZvLjdC3EqpXeOXPrG04hK6SGqY20yVN0UF5ZQtePfHM55Up56d
YZU3yMUoeCU8y5TufFYOTxrP5k9uBLqYEDQesfnwYSZxHha2/Z0lw5y19JnGSmS606G8yySEBDBm
qSXnS+/DeGs+EAiGaCZBdf0bpfy8VMtkNwMGKHCGN1ZxDgKVJByxtI+NShnSWce+VnHUFVGW5vSa
RehDdstVcE7N9/CDsFZHUushflSDTYPc36Jum1UP0HsOpkUBK2fLFmHzKlF688slmMgoCTa7Nj40
vhNaQdNCVGfTdzp4ve4eRa+JopTZsP03E2KcWVt6YS7rVYWpPTg2CPOhctfFrTPGZSCQPZ1e/KkL
yd6grflxfaG/oRc8sk9aXxvcttmDzymisHwprv2SPveNFDPgKBAlX/I8NjQDhIb9hlLJbQCoC7Bc
Zn4lrTBvg9atJOib5PCA8lch6PuG0+tcitSNfWVSHWC9heV8GPmT24lJw248pKdCXCKcoEFtIcMa
fmgOtAVIRFTgxvfMhVs2zxq48AdDakwfRGwe9wvPVDxL3wkQK5xFYzCpnEmvU1MWQOO1XPU9YkcR
A/XluJ/p5ubea9WDdCAgWdxnUMeASo73mGF55GbwQlv+JdL/Cem7IiMlb2o34xKOxt08BQnfk22i
RhZuH472d1ksaq5gbgUwr3ITpVXvtOD5J2w7t4GJ51XIeaiqrl5N/Y8JddGh9U47IzROuAnBT/bx
hyQFvCPxVzntFpG/iXxdSd7IYnDyPSx0L8rN9PBuTaP8P+10q922A4KhTS0DO70DQr7UZ/NYYc/6
/0i6A8Gm0irUZgmDh7QDYzC1TNULSMbe8nMe3pdIgu2qY+/5eldAQ9SnTLosJX1hm9S+gVMxlSgH
698MvQy0iW9/pdwkc/vFV+RWO5mUDKhFeRuKbz6CYlFnCcCJ87dVn4zZd3oOAzOXSOKvKArIkrvL
OS9QNC+R+bh/kTajDctgVyJJTueMU2QAzg0BDpGWTmGv21uNMTBD598Lns+CwQFjriCot+f6v40H
rOHzQpbmXlnth/LB/BgZxckUL0vUUnv9QP41sVGO79QjCE2EqDDht4wvIQQqnO4lnNfIt6eneGX8
wwgVdVRApDjAvJGzdbVeDEcwzpBL7DeB7eYn8brYYeC1ADjDsQmVQJh0c90C6za7liHRy6RYjiNe
Vq3GMXt2y1WYd3gkdU7YfQX4OirNWvwm1kdenaxvQvrsXgbnddma4G9hIrVQnpS4IKE6BrB1+aGn
rgQO062/C9Y1Ku8IQD4iZiP1kU6LEz/oFzNm1ht5nmE56p7nLSQauSkbzw7eevRnSuwUZKXvgbZD
Z+ecy0NbaYPWI6DEBEP9oN+bBgcdvPDIsLOupT+F2d5ib86S+o8WuXXU3hsheSL69Bz0hfomuttx
gqTPvMGQaydslalv1VqBbTIVNNc1J1YlgeNFf0ORr8vGrqqBJESeCIUYzPeltYCwbpUCR3COovR4
X8RyRPBFkCzRV8KEchPVsPnZwmTUbrPp2+d5gUYMZG/DYkblQUAw8btIu+/j5ULVFmdgJfRqzN2j
Pvk3pSns4H8iKucef9d5tdH58Lea6MYOKOH5DkOv8hKMYZCiohAnbt4HOIVavhoaSnPZ+YYgJ2RA
F/JeC0751zyHeHKaZuc8V/W3TrFFlum9V9ofe6AmJST2oQISIr14p7gYdlc3KeiFgAyeZ0fpBXjf
+L7+sbn5w9o+ceuCNaBV4rWtV+oucAoqEMSyJxoq4WPmmeNAjDq3AwMbdVld7hmaGcfVHnMGLWJj
eBWpO8Xt9ofNz2336YJPjw1JNGPhim8kfNOn5QxA9C+ARNsXDy++LYwG97j1ulu0fcEbJKRYTIfE
UM7+rZn8jgZUAQRDJSSICRxE0SLbQ9aItw3wqkjmp9gXxqevvrEd03oklZ6WrppzB37M/4e+sh4l
Ny+2g7SAGeXphEnN0TkobpoTVbSnk21oqwd584ZEFqsP3Ebk18/eBHj6YsTluXYCKsClnFU46jf9
Sl3fXyPlCxDPdCPn18NnvIkGoFYRK8S8vUe9hlmINv3PtzJrEEjbEUHs5MW74NJ23xfURQOxo3q5
YviaRqVTeGrt6VOhYYaFI/N7a7cKIuXZW398xwNNAYJ+g3m/+jIjM5ODntvaqOiRHZw+yG1jR4gQ
oBOEvCYBDXIZF8jtAMLEufGLSo4gawbz2HZ0rxW5MPCYDd8LSSgNuUTqb/Pz5nYfhZumES/xZzwJ
AjgsjdqOVP1INwZc/74Zz4kR2vJOhgY4+uBdEbLdDNP47XSr2jkyf14l7OuuDINb8bLDoXafQUwD
ChrY588/qpwx3J83oRzRwCat5Sg0H8SkhxSCfTqVNagmn2Fl9m2CYCnO6zmqYNW5REJ9j5gaUARS
a3ojo1ggTvsfiEbJtlTgm6ZyRM3R1Mjl8ot7kcxFDNeie6i2UK/kFSSzDgCPtrjS/m3uYJqoUyG3
d4h0wnVVWH4AVZJiA2TG9FgcOYWQe2N3oMO/mNBBTUT5pAnr7Hrlup87Hou2XehIsje014NXgh3V
kqq5+K9AeYutq1Gc4w45UKvlzBXA3vL/wfjMBtNT2pxLxenbbSH7+brtPNmZUXaaLyP9kv1aAZ/N
OPL63noQnKTTQ1iJEbCPB7t96UlaPffrUEGPJZ6j2pNdENeyD8QMAMyLHqgZW7IYPkESMjb1t/0Y
ptrhwMc4a6LG9Zql7Y9ryTUqhrn0deoLNW1pe1U75miZx3sJqWCJiZP+CiCDp7CSVRCUHDY9DEHG
58qW31r2SpdMdeB/1lToYukSkZsswOQM3rOlzZER3698yGDgfcURvimkEfB4cgMrl9Mho18O4s1z
LdVrdU+gxbfeSVRf6U9BhZ9AkKiD2aChr+tUr8+iM4If0udyaqsp5DVp1IhFNHi3KBcBqtNfWlxF
R3MGnSsNVExR/3gaqjcB03yMwgbiBTzaREvc4vRl8GrpXmyCjLyPU7qPFbWi7P6yiuG+7ki1Nhp8
7yfIkMwZ0N/BgmElnrnUqbn4A9DBILkYWOsDQFicrbCYKegHGSS5jc8o6P19GISSZjaoSx7kP0/B
dvRrCDR9Q3JVPz17UrhPtfIp73JlaeDD/Ddx00MGxQVZqieM0bqvqSsxGj3iXrFUfd7JCUdpw2dM
iAAuR8pR/8GGQKcq8X0vB54gE28f0HxLdLOmCDG8W252qyNWJNRvoJZfNwy8aZkvJtnBTu7tmz/4
beKleIO9Dr9SNnbShGINRTNl4YY2pc3h+IQ4kYQ3up7a/tG1iO7gcvQCDvSR3b0PnMU6bFkLXQdl
7RUVXNea+CbnItO0fSvvN+++IOqYXrprxe+SmEg2A4ZGgnKK+NM7mkP/TD8vDlTNOEy9vq4YrEUr
RhJfWR9f1FJs/fQQq3aYgxv0vskHvZqQpxR1lD9fOSbMJbFtQDWUj2Nc3mktrhSAM0+GfZiyCCMa
UhP63RoO3Phke2QxHRZuILuRLXCCG2JzponufRxd4bWfeTGQvUrFEzr+e+4P+d+So3e/KwGUkkSw
3oqHVnrvALyVRUeD3M6lkWLTIjs636Yc2bkBJUcDe6I2HNCuYsc6y2/PJEhCdWye4B9JVnj+bnWw
upg7Q1GXf5QdCOtMHjQeYscsi6dKF/FlMenLQcooArCtjG9NqtImDzI5UfJVmvWBhS+okhu5ge6V
IfzVDMfu1fwoTrC/8lveAEuH4XDMEnd2dwV8jEEb8WNHigQKKf6GKKD93AqLqwq025ECYcJF69/W
S5wQaeKABomlsS3Cnhs9WCEcoRW27Fmfn7+Flj8a5XLuoUnQo6Kdu3V0XGcjO3+mX5zM2ft1JlIG
9Vm33gRhqPva1r2PaXbgc9661hhbb1HcQudpgyRPbwiWFukCZMPonioEUUFI3su1c3rJv7KsEWFE
pwRGMpxKUmoEr1lUwK/XiRWb/8JpP/q24N8wQqtjynw8sGwiGgxdRfU2pv2HXL84xnOrRJ2F+MIF
8VB61cTBkfc9yznsChKkXeiCSxXBY0tXZJKbBUWFU657KbvnITdG2G8LADXVJNDBsp5ARyjM3AWB
EYTTYjVN2Qt0c8z0GZzu4fWyS3Gq/JirzLyFvSwFm67rCgac/eB9RRaxPj45bwzbnpEdtTPQzEeo
drWyG+pWWRIa1IufaeiSRJFocW9q3weikyX6qOqMT5HS0U76T9MV9rFN4HhqB4+5hnxtN1MFq6M1
K/XxUgtaiWkQ5E+kfEP6iWb7clAa+bLqses64bxAcp2UPLLu4bF46Avw0V8MZeaUFufnRMNcB9Ov
v0BHLhmMu5itrdajuSYH0nOdsdo2TMJ5ApnZLlPHgv9dxuU71PkGn91CjOdv9BJqwvBEeIfU5FXE
sYq+376Oi8Qn51mHQtBhRK8rB+NPAVj1Wb7YUaH4c6VwS0aXu1U9G/zuzAvCd8zjSqTHMKOlHJi0
FCOS3gLJwve3vX7dhR5y1oI1NH3cUzGw3/M+XCpfzrt0P9E4+Pkt8L1Ny1G/OU9b5sKYQDftoWE+
CiZe06I3ZxV5Sz1Emz9pKOIpezeV1DOSrEhFzQLiLUzuBTobZixWkSWa3cZ5CIDZuWS9TtTAnGba
zCLZ8xSfi4yfHRJqJIYbRLdjfjmfGaWFGVPdJa1vkHWasXmBX2KmglqsNF2/XN9BThsbaTesLlBk
L1tpC3yxegw0bc20zrbKxeiepxvfBy+b6Yc9q0TdX37VSc0pkW/SRfDaWYQt6yejPcU5CCLmqNR7
luk0PNNaCRlQjMDMeOYLJAjrRw4X044EAGtnsW4m/Cb1CYF/FF/d6LfcrNCXK058YZZ6AKe69jE3
znnIFHoKWqNJklQqSJryp5bNVDnPFXEF6RN75O0/PMrgm8ZXiD0CnOawPVwI8criyviE2WMd7VD9
qrhgDEzJEAYI5uPGWB3yPvVYqX73irrN16sQsPwk87V9hGwmWU0i1nOv4wNmotLqN5dZTYyPPhrh
m53IDBohploEQ7MiibO792g94tMCNfr8UXT7Dh3wseDYMFOOfXWSCVkQwaCCVbJ20XJ5gxx7/eRJ
hwQnyA4vtugkE5iMgCbN9dNlKjZq/CMVooSBQK+6yCVJFiY5uVwop6NTnr0bknCogmIdoZzZulh+
wimg8I5i1QhK5aluWd0NO/562CkwJbicdDkIccwlXk/U6e215RwXuw+8KmxuUqjvJgeVJhH2+EmY
ccgyx5PA+eeraMP9K/dupcutrJteu1GYFlU+29v6UNyVGBEvko33d3w8YQwSC0H+gTvOfxujeetH
E3m7C+UrjctIXCYXVAi6RhIMB+a2QH2S5LX3X3l28bk87N/A4bqUghXIZblLNYxEaxDtmBiQzl0j
vr8CSXLxiBWMXdPnMb1Mp96YapxW7YPcTCO1XGVXnaSn/73F+iR1EHIjQC6YqWotmtwNIDtkYQf9
3uU9hjtDCTNWd1gsCYwVuLpxMuwgJTrGwhssdL6khZooxfHSHg1/2aA0AGPZI8YOBaXWFtd+GVrc
g7+fqDiHCaL1kDSJv7bGrkwNvuVUqdHZD1rCWiouKvOXNWIUrmOPKlFvTWLNVwEQHovBCD4l46OB
ywPU3tvPqJNXD2oaBOYlMHxH0gH6RXyIi6IAqlIHGkI/XaI0oXG6uWi62HcGRIvje2v3u1q3/kJ/
VU5cgortN0uO0eOf+QdrrbiTipCct5ZAJdt6cssMAItuuwbE1dX+eR9xdOE3WPhx5QvUMLMhhYwB
N76axjxh5lKqAjqWnwk99R9/nXCmuVsd8wcxeR3Ci/jlvaYC5WLxNjLyHfRmuPPcMR5Yd8JxI25b
XyCkLFEFSZwgN/JqV+Jg+RDB7tnFl9ACLFvi+TjDedui8+eB7qQSoCvw4A1MiYiCE6ahi645+YFv
Kn6Wn9/YAvNVO9xcWSKAyODHKwbENbyrHLZjSg7dmmL6O9g+LCICgFRPz/ZWJMZUEGWe7BAx/yyw
B05WNGpkGwaaJHr4FK4HHbliwqhOf8uXgFgJGTK6PqZgtl0rF02U9ah0Nyc4lD8CpxIHi14vJmvP
j9il1o5nmq4Yz9xStu7qOpOCOluMQHMzINdUthd+OPC4vJ/kheR0Z99eJKniH37yM8c8jm9mDGAd
JoyUv9RZRqSRPKm1tOhqAQsJcTgW6IeM3aJJFFV88e9iI4F4lVRpji/xSVsC2tGd4GXvC2coQELf
KdeM9080O5sng+OVbdR+uqBAMPWZqbeZdq0UqSuQtRS0RCIvuRDgm2twmWIUZrjhGpNGK0iWw4Gn
NUOb7Y6EeyxEuuUr88S4HsVQcKgrdNdvILm+MEuzRYBgEDzDpV2bfbfKIgjFlNzhPd1TgyijzT4v
O3GC/3U3eReqP2xhrLUbWz+OxA/Tq0sc7Fjy04/rs5W3UEj/LJ8+k+HAWYUltdd6GD8FUfLdZnKt
DqxOHzC5SpCqk2G/tXQBtbltUllf5jzWGi7dZYkFdRw/KhOVft0EmbkrUaSJpjwYgJv3YKRegleL
FKM1mG1PT6F3miBePf3iOD3MCeZrY8z/3rdL/p4zE2dLTo8MZQb0mfaijaojzAvipDnLI+pmx+rD
3r11l7G/8nbiHTUGvzx2kkb2EwZhNmcjbltjyxvXaAUdPAo15iTIyTm34mYd8KUshmTq76JhIM3f
GruANc6BUXotygiwh70aL+inRrFPaiFbC6Mzg/WfmL/b1CXwpLKP4xPlxq5ss0HR6D5TQm/rF17g
N7vNdp2Lw9GB32UJOMrG/uvEAiqut+CFWhtnc7guaXgGCNzQIxi6xHgZgPccC8Tm5OhiI/H7DjLz
a23LqWPUA0j9+e4YVgHhrzj3HYSDnaVU26vqkU9ftW659KyUQiGodPlkMp+wDGJ7GlR5L2wCk1rf
M8IWUZVv/uOYQ1auib/ZsBXsCraZFSpaxoZ/VvPwljv9NIYdvYL++rBa7Vb6wHP4rRT6yAgg1rSo
gT/mn5L1FKqesO5Em6yPFo42BRH2RFtU8s5myfy4O0uHTGB1/CjsAleDntSHObDpj9a6LUGvRTrl
ZZhqWGJOHcVd4aq+yKvUMCkV5LvzOMKO0H0zYQLwMISMphw6F2yItnsVi6cjEmuPho6HadCutX21
5XTPtjziwm7aV3TV4ZMwVRtTVYxhHq5VFJUSQIHRDnGVeA0KIm/kowF4UKpKnxdt3yweNgk8LYaa
RtCs0SjRLHykaX6Z98XuO+wvsua7WfuB/MLZw8fWNsahA6XhkUm0p26eg9+DvQgyhO0L17A0PRXp
31aUlEF3buEK6ldqv2gNE++r4DTdbdOLFmBFBIxBg9DFLA+TbZpqNde1MgdinXOwlA8KtvFne8Nh
5vp/l3nnoSdKgJE4JwBHhWoEwsD+MRyg4CLoSAGKBbIqKJs61oCbQUF+C2J0W3oUupr3t1KLw7Yw
rChFmwggatdHVcrILJJyiMYGPRsyGo0JU2oJWuwnNzU6qrpCOiEgL+Z8DIFQ8S477nFaHGr25gO+
W7S6rsQH67HTLvyYTV0H7Zjl7cXSXso+wICKD0rk4UqruiM0cqCNm75uXgUblRsyxFCgJszJetjo
m+W4k8/FhRwWvJfAwhERyso5O/A8Iu7YkSt9q5ko4x+3zGpZPHDHiabEfl6ILFqaCE8sdaRuKFRi
OrmUSZU2VHFR9abuvU7xPcRj7jr2Jh/dD7TCdSOaCppY2nWrQZ5FovQCQhGMia2ge8hU3ynBSzoU
or3UVrplH3AVquz0mdsAODP/f3cM14BFn+moryzb2U/qmyhSpcvKQW8PEYRv81gboJpB7tOAJ55+
+3diIGqaHFtYuVBc17P4rH9FiUJ8SYTc6S5OLPlgokfwE9iBsZBPM20TnXQaPLVr4Y1+MdNnohaq
pb9PvNNraY+zHgz2d5PB7cgy0RzEFsKDxJVdG2YyhnZwVT0sG5Kd2ZmV5ztn0i1WJsGtCbBk53Z0
J2k9fhm1xNNPqJuEN7t9UhEGdnVyIkQ4YFMFKj9nXVbq/Bv2YVVOkGFdZirH1nwLI65UMYUoMmOX
FsURH2LqER3wtRN/nREnzOGfHjN2lIFVdskSe3d6z0c/Shi00WtNZnNxQvezsIQ6/ZQzprX1KIGK
W2cGY1rtZjwxPj/msQPYqSDfBOh6aJnwB5z7HEt5ulLxKa21SbTKv3Y75lFi8qfrIm+Gi5ZuSXsu
6/AoyUC8NVorKqsXlCvhKHMOlJmjaQzO0On+bidM/fwfUjewFvMwrpuPXSCHh3iBQ6/ULhyfk68L
GS2U9q4ZEfMyT0y4HSlTzTtkpL4Tt9aZ0yW9mesVA7Y6JOJQiavqHoR5iPdw8ZDSGfPag/XKPNmX
bvzyoRjHAb3Fz1cFQq9912hATWQzj3Bn3cWSa0sVEdx6AogTECngYQ5KszyfTgKCd2jScQHkPkzU
iI3f4c4WB7lNf7C360jjE9vkno8tkSMycFMYzDboxpWC/3JTzybMrVgtTwrtiZ9ZCISb7WQIqS1m
dd1dxUNUdODDIHZn7d7/zKhboKcXX0q7C1b0HTYyRWfkIofrhP2RrvNj5L37Sd0oe4L6wGxse6bl
0t6auHwdIUXBfmNyD9yAC5yLxyPmJ+QDMVUBJ8A0Zso8Zm2+z1GOGVz8bB62E9cLdQsYL/xBVOmq
Zij/s8UIp2S0up7VSzBm+3lAY+CQLChwQkxVGS/yJ9FnGJHNeWx8+AUdlCvJRQppalUAl7kPRZsn
N8ePOfkgT4y1Rx9A2fwqapGCc2jJGQybxFN+VwQ5U/uo0cL6qYBZ4UpLzWgeLp8H/I5cv1tVuap/
33aSYUOqvw5HjYiI/Myor81FYeq+XXkYMLrzyn85K4K4ENWDWmyWXkXdlk2Wz7ECZ1zTEE/eE7v/
G+w8UWkpGwRQ3VnTNoYEaNYU4L/OIEHn1uBGavs6UX4t5RbQ17lxxzfURBGrzfAD3a1R67GAuJyT
LF3ND9LTbJ5yCddYPJn+RbW1th7DVDJXMpIY8Efrqr6A1NxqSQp/VqmUv3wG2y7mU0R/snZamrWa
P5goK6w9JbttfrcNqvFluINnsPUipagQLCGh7F49mS+3OG3nPpphkBPHm2i2AjbxuwyUfVOa09w0
GLPJCk9JvnGWgU+ge5IXS+MCRvN3pqUBHG05L91Ho/sh9t8uta71u0NDoef7Eq0ruF3DfJI07NWO
Pmb5Ri+HtbsR4k+YBjbT/Cz5OQOe5dTXOoJg6mOz254Dh5LzdkmibKge56wSdPQYbF6F9LxixCb3
vWkbX5/q+iEoZ3WSMKJbL5wV5WbIhqyzqV7VY59dvtkMBHzUsyMo44e+osBYEXgDDJSH3aHy3kLn
KS8THZ0m8d5yc8/V6+bRBrxwmIdcTrBvZydU61gkMaVqYQJpPqjxbatve3khzx/Z8RrYP0VE1eP9
vLOLbbw2z8mIVwsGDo5DzBh6lXhRsXz78+0GS/hLaQfKqi5R9AWS0jBFfFemH/O1iehSSe8DxFs6
pTQXv2qcCYBMP0ib0dtGeaCh2EmSSTPzsPa+kU5emszEaunSIXJFSH1cLh1Xk6p/oGBUJk7Xmf4z
R9dKLiYbNTOjHjwDCMaOTRfoGM429Qdx99eflnqB4y3dff965+K19DOMNU3q5LUt+u10Kjv86KLV
FWZDHmjIW/xWHaPcrmSJAMK7k2zdQ2lzrn59XZOPQTJY6vDmmW0p9/djwSOV+0t+1MZiZmK4vfks
/Cr69Ih4aVqdtJE4j7egKTT8MlQF8kt+Mn/TVQG3XWJWxcEQWGuvjD22mbnZkjkuMmvXQX9aEGG/
yaHPaQBAYn8d5m+i6J336P3AaF5bWVLgZtYue59Q7AYqoitB2IyJU5oBHenPFE39fpJSrambA57L
6HRkDPMyQ6zld8XP+ox0bWL5UUf16lCcyyKEdnKFpGLHhRCePdPUbDIUXfK0jCpgKIT0otnQvXHM
rC7mHTwqqnvuXNP/KIb0vlV0hjOFy4qFmeXydHEmIQrkhHFG5GPfelRFPT9wNGUJWrsJCIOKWdGS
sJbN2Is7hqIRLUISVW9IgsIwQ/5cTnMj33RIJIo7VF/4Ex0cX/4U6VicOnoNv2Wfv2RFxvk6Rcrw
p9y0BBcugTCd3RwFohnqG7os1CsMoNVOYzB+GLLb1pjCqAyceggi1ry1IatbJ5wakDOcgmlF3vVu
mM+dafHnbdwJvT5qIllDsY4pNHFqCpzYShsHaU2ieknmqEMl4aKIwaynFEENHZM/F9p43zCt1Ifi
p24b2d2xMnqixAq1OizNz4bcwZIGcyTICkO4vHoXvkZQG8C+AxIvtcqtEOCqiBgzGKOMEKGqbiPp
qUrSF6xpYPEeH7JyBCN2r6Ysb6WGiZE4BUAtFpxDWS73ZM1fostsrc5HHnFBGqutOqluz4i4jf8R
hMfrxCtSljASdeP9N8Edflf4iuHqmnlwh6wCWFw1WoGdbozAdWWhw2yRwmvyYc4qPNPn4QO3IL2J
uZs5WMu6khAovQquyycVekjZ7mgfaoieO6R373XwKPZR/LJWzo9gMrtGAuu+pA8OhPpmh804F4CB
aEA/woOEYAitpCMJz8kiha6InXYbBewNLyZ7GoAh5JVx0THfKNxcubUQ9HksEHT7C2BqnAQF6n/C
UZNLv3mmiSIU3apmAHH6gvh1XwLpS0aS+/WwZoaKPqr/exPg6b3STxwaHXWyKSNIFEig5PCkl6cD
zwPWzjH89WelUNQZiXHxEwY93CMD1JvkSPcP7mAKHcTGO0v3J/OrL5k6eNgJKS/7pTvgY8GZH/fD
JrFVZbJpx1GLcaS+Y+jdzIjx2ZYgrOZ0a1KE6vYcml5j/8u9WNZCdlyqmCpqC9Bxf2gF7gHod4vt
uasvlkBLQ5yW/s1MqycUBQhwBPhiWzVOwElr5a7ucO1yUV8Zef1fb+VFSuIie8f+xNrPKp6p96h8
m1Yz6FoEmt+BLF4CQw2w0JiLZnWFPwxt5cJZXbTyjhTEg7iuCO6e4TdimECNHAf+hY0807R32jrU
muQ2RdGyYth24s8HLmFojNbvPlt6b73HKaAIYXRYiZR+JIfSPxd3M51bBOiRumSUUURlEUfcUwmM
QHRje+eIPm92YLRqtLBJ+TRJ+Zk2NHHlZsE9aUZVrM3rwkkPg1r3dwdd9w2neuamTEHSSEjRquby
JJCuIzGvBlT7VoaSAC6KuPKw1cCJKfISUOIFyOTEB4vMI99SqmLg4azLSamXH2GWiabiWx7QXfaG
Zv4JXJLRohofzUnAar2Eir/1w1khYCOZ437rV4OV4wJByagLIefLcXF99k7QYWUGaU4754zzsp1a
tR0c83JeToAZ5oyFUE+8kep0ZK1Azc3/Du/tfSqskqatpRDDAaTF45hXAoeP8hPBJak72IAYurns
8f+cN6pgPRoicLxeefrUyI3Cl4GQYYKvl4J0+bdTE7ncC3QNHsLQuFQ73SBEIC+U5mZ0iCw1LOwD
QG0Mxoa8iKqsFivmeyQKSv6IphoPZIwIgxq26/+MMY+wCHA/CwDrZdDtPBznplSs0CaXE6ecYXAD
aGmROtMUk0qeLCLz3JDtO6vVYj7FH6dfbvaQp6Ge+qgxrwqEVuXES258LgXNK5cu9W04agzzT8ht
R0wQeQtHPFhbL2JJZrXcg6nVfL3BuSLbj+UrUYBQw+3cB86I3TqZeOww75ztAuw1621WG4r1vTCz
NBVWdMi3RJ6IsEtVVI94mfNs+KZj9xVHUH6yNJlvqCAl5VrlF0GmPEXBRwVgqwZhj31VrRwbXJR5
jULYVGKsK5uufRsd6hQTipGuE3bUOXdRAQLKXQEv5kVVmcY5oVZCd54wMRjQAUHupVxAjQ1EoBzX
CE1nY9A5mPypy7baT+fuVpRH+zQ0JV4PGdrMQqoUQHZ8SwB1+6G7K04GM9+wQ6iqgUaY3xCAMQuD
CzUlmn1SQA8jqwchjWpf10aV62IrOMZ6HCDXvVjIFg887RKEwEeO51xeL1r8XU36fH40W2CY6tfR
EMQtzOOhlxLoxyDZbuEGLqXHm8phGjuKz273aX1t8B+bK4f/eONr6YSrXm22/3B2s6sEBav/cQ92
kolbIjrVm08YN7i+3CPytn9yExn3USBn82d6t8lJcDtV/PVHJVCMyeyRRkRrPyP0WXldkkbRGhhG
haf3fLwALzkQRaHHna67ai0FWYH8h6xgttmHeyO3vjQYN8if0GibQeBx/34OSxQI4bRL1nTkXZXO
CyuXCZNBxAWMdIuXv9b1QcsVbksofcbBCt+K86wK1q7VuihBlqocOcbTO5RtuOYs5xMcnooafx+k
iSGfx9Uhyjr1V8vjCY0E5VmEht5O0OiM/D0bwnroPx2Z0fq+6j6xC4K3iLwVDNaZoJFYSSmxsZfA
uMonScmCjwDWoem3mcNDmFtqmYGcLcTIQ8lm1IGSHiPY2PXB8KCsAZRa/cG1j8DM7Dff/jZZ6RBK
5UcgdlpBn/Dw/8XakrHeOL0STonP8fZiFFWwNo8MFyHSG/5dipp/vt2/xhbuvLywTCUn0fpB+EWK
oBa3qhp9la1uprDA+F+0QemeMZUJQX0EwJCK0ppOsyXPT7ob2XDTORuzQX1nCgysmheAANSUc70R
Zi13PNpHfuUkfxAQNQUhUg5Uc7lQNJmnh9MiPX+9IuoJF6YOQ69ryXQZ57MiX10FUQway8/pFvtX
HyxHky4PjZms67F/AMWy22Hg41MmFii6ZCAKogxHnTKU8bHWUEPzdeSoq89MmLZcrwBXa6UkdOSo
kvHMzcMv+ffOoptUvb72hZ6JvE+iJsvtcEO+BSRT4637EcOO6NhFrGnsiwb/8cLtYSnszC5p0HW9
ZiZR8suM6lOSpDfoppqxmS4uQn+VAJ6jV51Yo5gky9G4PGm6yqIrw1d7NDalfJoY4U0WJWTytXt6
/ZQo4KEumrLoKtV5MyLj527cAvCJwaVff/B5Z/C1T0x5hvMpOsQUZdtxBLYVclQxu5eq7Xg6fZdT
COCq87MbNULtBhwPCRfbwEPmb9Mnf003QALBK7dTDgT9yQoJkzCSEbW3w6HUbrcciacaf6IaZyU8
i98u8sNjbgGWm4y8DwyD2Dx602rbmetAGVtNf7Ef1xUynjtG0N5WT7DFYlGrwqHDbxVX/qvUgsSY
xFEPVy5MjESpCCIsM0rZlPPupCNsc1rWMXik2ypotyctZiTvWVTgE9iYy/Wb1yu8DP7uBsW2029n
03jRxNXayo9zEQLrqHcUicJtxgKjy1wuRDvGj0R279x7HQPWp9glpj7g2Ez6wAaP4bUDr5W/kEpz
XihFxu7qmlJN1grxAmEmO+JCdh9XbFueFiORyT2b1kkPE90Q8cjablOBz1zrR2gogMgrw9fRMt8t
weUae6WOdTzM4JpXQbHNotHB8FEbi1rtvsqemB6xlwVNV8RwyMwoqCrulijoA/m7vk3cKoY6Vqyl
8h3RnjU5GRXDGKWVBz2KLk4Y2yzIN+poA28T0jVdA+3RX9/2dJIJ8CPd6DQj1RAi+fllkuI9Vz/D
/ZKLUSy9OWLbQ2q6COsb0NNMkGxoivpMYQ/mjTOIM08RvMPxDYdLL/Ngff20D/X2Il6Q6NcyH0OC
eLu+Yjdd7oN7j7SXvePU9FSvCopd5kq1fHMfyDrxoh95L1T2RpBmpvFRsvPqyDEeDncPyj/8o65H
7zH9YHPtA0alLHYtwfrDsVHu0YuovK1dKeaHmjDnBQ//4oURc36Y/MEzXpFnndWAa5Y2tSsB6II5
YQcicMbtXqp3nRLEYN+AHttpWK4s809EGW2w7nVMXsQmiPQQdAnsqPKmZU8rYan1U77V5AbTNkvF
7IhFSMLj189qtq+5zvKovUo48nmUNF4fFzHrt8v+PNAbslAtrcZ9ko5KL+Y35yHdzfsQpRF+5yg1
B0LyCyWhVtoPVWWLIIA0LUp5WgO4hv8MBstd/fQDOgaJLO3EItNWJn/eUM+qWPAKVUnrX9vH4M2B
KYOatuU1qklJsS94OsjahkMOUX/ch5JCMs3zgZTEwwaF8FjiygMzhpZh7vuvLsiPedzTNNMeCghr
7XSg70sP8yE+qbx3okjlENe7aTVOcterGxIJQBUGUyGvuXWzcUs+xxpFN3bfhuxM6x81DLIzBUJI
WIBsjR7YtldKgfLQEhiNqL4eapErfKVdXpxkZlqJPPhP6xBIJToZCcCTfpb/7/yDLwc6z55CnWy5
RHpg18xrSDNiwECvuQtjWpYOHAqSrguGAeyf4grNr7X6WmoETgpip4SsrMhB81cN24tuM+HYHuYV
SWf4fgQu30sOZwCYooO+muEw6RxsfZMyDicNSq4Kv0/SgPKha/6IsnSbpY6ygRx8xm7wjsPFg+p2
AKSkKkaKdrMcD6XiSip/M/EbTh8xLGz9MO9VqXOae7LJv520abQtQanscMwv27wj3GsMVOY086Uh
l8eTR7NTkQq78OYpxBblfDrpMYB+g/2aadK3RnSAolxIY+9ak1aIph7hdcVjEs97MC6BtS6DbBtP
l/M3HK4I35zH+ZBO8Hd7mcBAlVWN8ttmt9RbvOAquu7GVrP7c/mxJrfwOAhAnAinFY+w1ZeyE4mP
bla1e++NU78fcWOyV3Sh8HWqfZ600M0s3GqHvL3uWbEdt7ZxLvPnojfeqd5Cajwa79Bpgm3YlExu
p2ABA+q9NOVPK6jHz3Gr3nn5aeP8MES+dLuTM8PNfGeWGAi5a8sYuRqDKjHv7YGED+vMnqDGroAK
MS9sPT3b3XtB9DymsDyLLA2Qu3YYkyL/uTFrIqjM6fzObtntC7gogoaRX17Efa0od3+9RkTs87sk
wAodEwWOcrbQZdQ6no9j/S4oBfyw/ZMxLCVpzem72Tf9EPG8hl+hA8u5l3d51Nl1uLSamu0cZ/82
F9PgFMXfsE4GIqlY8+DzjMJ47Cym8sRcqrO5B0CPvC2h+jpywBEmPrR0L9BOw4iuiKVGWsRLkvBS
KPNTxQLcK9xaCFvERFVaNro3AQyX9lysNxS3a5aQZXBfmiPxttEFFhcETouZgYcntEImL9WZg5jc
KL9KXxZNcltLRESPTF2APvEYFiO4uqQ8Bdfvr4of1sVuQiU+DgbX7uWPG2D/D9RzsUkisCxaCuvs
jyNcg9d5bkQzyTb0jPHoq4fRYmVa1cVksaee8Wtc4QiNoulooiSM4yxeNFqLnJ8H8EuoQQIIpR4G
ykIruA7rvwtKMAnvu6Fpj7I7y13ynF6aWD2NKzxYW09NzGJNouVS/l1VzrOFx6lwb6eeC4nDatVz
DDcNeV2gKWyxXksURZI+HIJeK8PoFIv4jFwfsDv4nKBTBfI5/4OzR0uQst5Y/xDxXpUlpMWKQlO0
O3XPpurlc1JZay8m/9j+7xAHXgmRRF0OIh0oKz9bl/6yWaz9+xkWxny70WChvvhpIu3wulQndNL+
E4bPebqOML2DtCgSwyZE6JOYYXlN1YI2xu4wqSxDluS1mSAQ8tkkeZAIjjLU023vXGdyxfR8vVIH
GVjGCT3x/aQu6/WGSZLBJJNouZaRX2NI0bn5YwSawu0v2MLMJz4xBs85KFCvduUfyV4Qti33suSD
nNsjm3R+vJ2KQtR4Z1d8kqLYNGjcH5wXLy/zVZP38c0YtYtBdxA1yguOix78t0JSrkHxfsw5G6Yp
YgbIWi1PKIE6sUchZfBwthAscl/ZFoxqhP+ZaddjQfQCPtYmNdxERYt+s0MOv9IXlVJg6J1W3ZXv
PL6ab1R/3TKWC2fIeIv/ewhwd4TTdx/ehOzz1NMy//wbCBr4xCL4IW0HnoOXgUwLtDv/0Hj3VLZn
J+si1WCa6tOMPBeN9/sjstsE7otTFYdh/dxawmkbCmpq0/CYWBTQK/qTbBLbeLPCmpc8kKVMkT5T
9cx/mROmmtxd2OhGsSxjtzR0ij0v2Gz/cWMWMaeHSTBqAuvb50uppnoIxjLFKCl2T0W04bJZNbGZ
I4sp9iD+13vYQupqr2cV8N4RZiX7I3bUd3fCrmMers0y1sgzvyNWPsyWUwWsKnwa7AlBI40a7GFN
pCEIWfQBiqk9G8ig4cIf+pRS4sE+uO8Cai+z7gLC5OI9N9Dc9cIvgdZJPHfMNj6RSm7MKBEXmOr3
c4+3c/CL8kjyypMONaP4ZwNukH1ZMZ1PgYfcmqHFG0u5YEP0A08zvAVgdIuQ/3jgjVXD83jVzOHZ
Qyr1h4GASeNsZiytrnvg5FZFqby++kN4r6Q6UMny+WQ2JLTU7tnlkollF2izT+Gu4dgmfKhMICDM
+g7vC0w5wytOWfDrVx1U9Tvw8FX69slWW8TxvncJSwnOQN2JVKLeqNS4s/Wh6IsBsCIvLqO2ybWf
LmcwBeGZQ5rAEosyq8A8wWaQOW6n1tQNG41pOSWXWAJS5AS/nnnU7Y/AYCqTrFRxFiIgHeLCcZFp
tPi0kIEOdBP541C0S+tl39Mxx4QPNoOm+uOCFQU4AsSUx9qry4N+QPvTBddEei/uN9m1sD2cfyMZ
Si5nJaAuzq8qDrfMKY0hwGDF/mPtr45urb8+AOOsQV/y3gBg5OCisGJiqMYI8NcnRb17qv9/fsGc
YKx/SYOZ5+kt99fpPv7LZgiburn/6DCI/nBRP5nlbJdjtIJ/OpE98XpvpgAVWsI4fGtBrgz11YAk
GPlMqdn6uuG4u6TjCH+/RA9CQUhm3HprYOfh4B4TnROqYdnDjjaB0go2mewvjS60Ki36iihHmKBA
6rHh0gaUTgWUJYx4uqm8cIz71IhvRdqb+uRnXdehx3QzntnM19pDwUlzBNVfYLdToMD/SwpsGdlh
w6+gc3ksXDfQhHn8RhQB+rIw66NJOZEU7vVZ1qCG1qTfOvyK+eK7DN9Z2Q4z/HKpyEEbOGtFEzHM
FMXQooM1hJ+rkMaRH/aK/lKu/6ZSLV3DeMZ+T5q+/slH/Wbddob3s5JeYdcg4hY4WX8MZKdbK/Yp
UjTPxPvxN6ZlK/aK7Srxv8Yqc1HoIEjuy65PA/aMokaFtUfgcTupfyXLcMx5A+5jWOmRWppbFmTH
tPE8DnoVb7tcuMkC0GCPjEVF4qUgKMmvmqXFDrYvXSYvtChJl/E/CbbW2nPDPh8436bdp+5D802D
fkr3nZVce6JweQOyYh6NQ9wlwZos5LqWD/xMogVq36or6YtCIAHb6qdhn2pAiIEOxQJsCufNAue3
2Cta7G1ckaFAJl5zFl/TUoLLQBS0gc3PE9m7h7yxZJoQWwrmGVx/xlI6gc4J9b0/z3wJxgkFMO/m
AKeHnsSnPW7Zh1gv/6oBqH6pbjoq2Fo5RU95vYwT9OMGPa25ZC2oR8ZR+Zw5+jPX56NSBmCELvVG
oPMO9+U+cT/CL/hYYDdvEI6NQsw5Jzx2LGXjkpBEwpNhDrt4KeuGGEIZ9gEbrSZMbN9vzX5jmUMz
TL9VaqI9ySG5an9K2l0DtbJ/whf4rcTnnD8Tqpt3AQmChzBiJP55FvP9SJAC2QSiG1iCWcU5rSif
RmaiQ8Ix3ayA7raXHvH9vdY/MGDC0vbF+07JlGqqOZAXW2dqoNG74rKAkUZhWwAwt0xqfMdsSRO6
k17HLY5I26amc6LRvkwubr4K7TUjLb7lLOG66dBSaJNgoFJXPt4vewAda2Apak9QC3aj4VN4+aKw
/ME2fa165cjOTcXd7aWrTowZ5nekKmFjZHLxfhmIcJcfJJrCc0IzZBKeEh2TJ29aInkb85evmmKl
Tf6cX8Zp2TeZVPw147KCprN7tERTWvRKR+wOON60O3r0mlGTiI/4zBJ8ubAQUHsg22woeRaIM8rM
/ZSSQui3eXzGjy4GxDLddwhNXNFxKxv7PSvDg/tdh4G8j418NV04T3KnZyf+qJQwMsui1QatQ9J2
GcwUhpMeLyCMMD+n9kZ5AHCYQ/vBEtb55vPWkNXZzj8ukdY8zjVC1ducuQYBsSHTI3okx3l8hofL
mLLkDPUiUC1vkWdZIOXYSwFVAKTHHdmQd5ge30FpSKoU++epqT+YQAAmaUaMGzj/iHWeBAEnydzw
5Qx5QygmK79BgbHs0dE5+L9E25b5lqsZNm+t6SLKJ52jLUrNUO3+4xt2siTrO8gaDrOJViyuNaCk
3nim7amZ3mmRlpIynd2ekFCr4/14F7S2oVgk53akaphgL6TlDBjbafSpOUcpctN7IxeVs5MV8Km8
uuhTlTv13q6oqTuOnJs8bYZZhQBfN2B7EGR7cRPCphSv6Vj42a7ECqNpLkpyApLVgCdHEe0HUGA2
4a9oW+0Jy5R4ffZ7mAwtv1If30yVzOdSDl5DYBKZAmc7//5RSx7+Wr1ia3Zz8KZTQ6zEcyWJoBja
sOeU59tgJok487KDgPpIUcgwTU6JfgxYSzW1uKMvlDMXancblqQXlr6pTo1Vxa6nOOW3gZSaMXnH
nM35w59QpUbACUb0RZVOU71TucQZ4wa5v/Z3FdraVqmo/MaMWVS9afc6/R9tSF/pMC900KsW6g/j
povBSTJx4qla2LWWgK5t1XTPyvxOI39VX3whcd4E5xEBPkmYG1wQluJzJneR6bkrx4ZrZ/r/s8o5
hd5GectW10NbTgVBZXkVmGNwTsREBkewFGBL3kbwnyx7EPOW6mnWHUSQghCVLmSQXGIdR2SqOoRi
wVFJZDHnY08ZVqGK5deE9Zhvugki327mzsQy4T/3HE2Miz6l8WhbLWZ/ZzYrUaf8gPK0YFa5Xb82
QN/barFEjxGH+2YDS0NMdRb8aczZdy74XYMRyXkEUZXOTEFmltnfhWchw7Lu/8soKfijV3HGBZQa
LqaAmslqUo1N0rqQvjuDxlCqYg27hS1b5JpKac18NFKgWO2wBk8ejYQOZqIAMrn5MyH6kX2hQ8PQ
wikjZuu6JuhBAle45Z/fi6b8MvL1vnARubuO0iwU3v4RKgYS9PPgY22wt2Sp5mbpB0R+AEegs68p
2ZG0+2KnvttfvA3bNg/UyXNiic22VAEGVeO9gcPWcIK6tzCejdwNOy5P0YfwTeRx/9/Z2G7jYNuo
+FZhaZUFY8hBwSuFnycB2SIXbZx+PvXbU2MY9ez3fOg7YeyHYcs754L5Ej7dcK/JouH8ocJxP/Af
dE0X/ZOH0eGb52IW7nfeuvZIJW4PIAw55zXntOeyubK8IpOiP4bLvYl0zZM3i2qkhNKvIGXUfLwk
17LFQReklXdA6UZKNubA0LFShRxTzTwXvGISQFtAUXb06aVh2J1jpK8r7P1vvHyotRk1t2aC8jHW
81dAQTezf83/l3nUo6El1d0Y84Hox/TuNRjwho3BMPPSRtNZvOwTEhvOEzbpNdIOhpoiCfRLKUAF
sbQiMc4/8q5H35HbvyJUA2RBqJO8QzzASMIXQkHbx5Lcy/uH4veK2w1iEkM69BJo3+VFdustUADo
wNAT2EEqy/JOSv1hMSF7KlFHG0+tfgZcrqvjSC3VM2qkEyW/6xuaYg0jJnSUJENE/0L/t76C1D6E
2oRal1Ju1wUGc/7rOOwDvnwqVFGRDB0DtplfcCiJ3VdA7w71kLOGcXq6Y+5MP/FjXdXn8+TNNSh2
5byakMgg+WgS23h08OVOSCqHCqeBBvmv8/doaZM0hH+0S1OU+3ESQaM7zm8YGNRY/H41DqSf7VLc
2hn1gnxYrSIoFIMW2yEs2fd38sKYZSrp1bhHU+1RARj47SbduDjCgBsKWrO5XOfE0AC0BE4Je7eu
xWREqPuda3KyshEkwWG1yh2JRjl4pkEeyFS2A87dZSA+1OvdrxgJIuVFlYIwMcY/pO/hhEPzBEJS
0TaRFT55TWBZzNbWZ88dJFZBu1hzRx27hjpFII6js4s/C30vBwjgTqAVpu531snaIJxvuC3aKM1B
EqfUA+bHNr6VkBF72AFNCXt5EsiOIJ1rCqBWOtzo3UkEU+hhcCTb2m1woKqv6alDDZiA3R8rxiMI
Zpqtg+GV9Rf1j0mFJtWHhtwqoEZlDxvStZJXeza1KUsDelZhGWmbQ5e3LCi12MBzgEmQWkk/yLU0
5uAJE8nf3NbdVmrunIo/dC9xg642k6dvF+9JGraOf3K8i6TVbxlMlNb4x3+JeqshO5o/e33qs9ch
gKiptedrtSHBWBUWH6TzqKDfWexT1K+8zJ7DwbzuViXolT9oQETnPqK6oHB1zM39DQXcOR89blas
YpHSBmjC/qQ666E38uDa3PyaS3gTpZegqkHBHLN3d0E9AZaR/PV+YpSpXTrtoKAEphjAAP/YnLhm
PEyCYWDsHV67i1f+l+SHreaDkE/d3tmJYKjER8ExGt0lhu3X6wPbiLujY9CkylJ5/GP49468j5fO
WvsFmePu0CM6Qh6H8OV1jPW8lwlvRPpaT+GT2UcUnUMmM5tF0ix4Z6+n8uTsJg1aVaiSKCre+qg2
iDkgYkhgQ/jrUbkiNqExK5HeROfDk3Kr1O5gV5IX1+6U7kXZDL/KkPmaJGBipbAOyMSaxp40iZ09
pdYsALEX1aEA8Srpa9VvYwYeloj/SgCW+YOM1/ZiUzZ6qnlrJWMk6iOH6tgSoH+rwP+LnWVRKir5
GBI3dh70DJyFWO+rUkHsLy4ddUYN37UoI6Xg0pZHLluMOO6v+SmqxMAstWDpue5ATR6hQPJZ5mBE
S0W9/gqAFE7RHznwQR2z1leS0OQ+9Y5Ut7jb6VSc4bePXKmsIqTULwB8GTZUc2LUIC2OQxLXJYR0
mOUOgyU2YPRUdZzF1DgTr9uLfT822Gx3BgIguPilzB40Qo1Lf+XW2f8v3EXpp7RM55axpw+Gi/NP
eMj6ArNTMpwDlieulU9N1fXOXdp+MB3dfvKFm644+RloIIu3oC4KFToLi4qZN+mhPRCuI5rose4X
2doeNOjSnepRzIXB3ZSAaMrwLMbuai2+aTx/h6zZgaBgPM5Fhg3MIlXqB1f1J+ylxjlLCb9aIhys
SFVHFVS6ckyncJM5R45aLd509XKWAjUdIWdivEsjGdy8L/nUo8z5xBZOZ/VOHN9EjsKvkGBTxOzO
NegPmbVX2ZNIv/FmFbqPnuPGDIAMd4TH01Gc3/zDNPD+xtG2C0CjBzNHWHtWYOeyRljnX2QL7F8z
QVUdOWzu0PRLK1Y81t9HSORinY5WHL7a2cU97YobcyU9GOEhahYdybSCQPz+H9toHOQWEsydTXA7
+RMOC075qmllBrijINjV09h00CHzILV54DOASYHvgUPejOJMWHULpJTmsINO124ajCwcs80bvpRL
9Az4RTKyqUa17Vxa2AV2q6e8EEQ4Syuoxr/P4CrN7wlYffrj136svw/qaNBrDaa67YSwQv5WCwvS
ZIbmPw6WPaqgVxde+ufKmbrMsouZkAYJ036WQJ1onolknPdC7yNxTQLUdM5EKBnPeWibT+Bw5Cd9
sTU0FbIZvpg/ZLhOCT0LFeJ6IMoYg0mP35TyYTXy9mHetAZBbvXaDbm0Bxe1zs7FJe69hKxkJEsu
zU4RnUgZArnhgvuZ8oYmtROsfZQEd3XQ2QyzNMbahnCV1eYj+CmJw9OfREESXHQ3yYQ3jMzySnbn
u6/qWVH3TuFMxMjAOD6KCjGJXUPNo/9zOwq+GassmiYNUNxBy0yWRwXZOvuPV5Gx7VCmjocknlBP
dqP2GvABvVg8jGxFtz+yDGpacD2IA0MyEnG7+pyd4ajUHWm0PNZnrhYPUAI0ijEaUIwb1RTfqW0N
lJzJgteI9Th8AlrDzlIwaBUHNSs9Cg3jQDUhFoaMIuz3XNxKhwNGkBvNu4xnrpnfw5jUUNep6yTF
gS8vlv23Ta0CYDmFo3oKqy/dmDnJhrQjHMBWh9eInX6nAa98ZB+RtMLcOtaO0WJNBkYJadgF52X1
SHzfiwin+YDIUyienBvMp6Stl724Hp/QITOXit0yqetv/DBQ8WhU+UzSobZe1eCyAFBG9IuDc6Gx
GlTt8uFmWeZfF/bcznlLDs9FdRhYfL4jd4/JZfc3kOYtvdFCeyBeDoEdQcAr5cnJqjWrWcA8Z7fG
ijjhyU9OHCe3uFS0hDmwviQUfD7q/JDyx3WXEn3mHKbzkQG4UKJuOj9UclrnuktnegUANnpnqx5i
LjYI2LdH1uA+n5FrNCjl2oo32kIBoCTcTNuUPdvnMLisL0jOauQoMbM3gcd0THXBwUSIhLnmXxKX
+xXx+Xk0pAcu8O2QAFtvYBCpQ2+tp1vWNdWmbknMJmx74kHlV1WIdflBxrbqerHK+HSHPPvoDRsN
4dW0P+c0wzZ9CBsDnNfqi610L9JQ4xEhnynY3yFcGumDumrFnvhUCQb+ZPp9IaLru9Z8jZka1aLJ
+BRTn3C5MXgYvbl9X5Kfa7whCeOhvTVdTVrgN7tfkJ1Sv0K73q19pPEmosXu/1QACjpubaPeLTXH
qu/BmZGe08Xdqf+8s3vAkOgQyfZp/9npXSRKcZNAuPflGKaGi73ofi9OsTtcFaYPBtERs0On65sM
QkW6zlbqj5oiajdKiiMFSXF+lwzqkc3EiKvCe0su0afmvqyXbfbnzBZx+kcWl+gMOo/umQH8pp+9
4c907Fjc2ZqACK17Zku4+h2+/mqiYDYzmueO4SyWYgOkv+oX620wC8X4w5OzzIuIc/n1hZwa7D1V
ync6EawL20nJzLoh/sS2mCN6Lh8oYUji2IyIZ5ny8ZRhydf7a4RvPwII2gZi+4g9V+QG/LmR6VNv
20Z1AOu+sgyYT90v8JFEXlRkzUrg3hxvf3/g8y2h91phGbrqBEbpnJi6dGVpNvSbwJNBqEJ9qFbA
94oAaX4kYi+ylny7ALXY7npqfltwbtboYx3xozmnfvLjq5nAEZOR+KXbV5+k1iYWm8b2YnqBcWEv
YZMyAv7UDXWSPBHZWgl1eCMt3BDauw2TkJrfi0qgY5wdGQWnAt7b+dtZDAlJ530wVKAqj3Odh/hd
eVj3mTu3FpuMaoGHa7sHrOiVBFzKvIv9FPJUvNavqtxttJME6+tj06/82RRAcXIhqhAnjlbxAxN9
SWPAZ1ewVttoHOgV9s36UHeThJewPvKZrvwfPqDemVNudhanPkSvn/z0j0cuDIHt9vkRrRLDyhg+
GT8YB8etipgBMPDNP6EGLc/bkN8bJj1MdpnzjJfY4qGa4gOvRZehsCubtHcP4UyMzqchhQanlcl2
b3M0vyZiXT6HDNZqtcGpq95WdtFB+vEnrMeAHZ0yPZM9mZ2qcUwr7eCjyQxUu/hKkSxbmS6MgZui
2RAMugUdb1L/LOGoxTgA1nLvLyCJ2TLdzQpaq0tWUluKOXQT/LdFy6o4pMIjnMNM7mCBIPJn+r4o
RLLcrhSGe8iOnIQbJcnav3L0oGu6A3Q2eKPDaqOj1Kw4naI53qJ80E8KxRa7qgY8Mn3NfQhsaGtp
gWruHQ6Y4S+1dWdER9f2G6g64Awfjs5r886O5S0AcfLpAwU27r7OGIWRMVfgHkQGz+9g+EVHEJox
hOP3sA/MhDFsVTVB3JgaW/QPEalo8BIy5uyifmna6GIsLJEkYLAUf+z5FaQgmEKgf+xEBUKzJZvS
vqEXFwCprxaqUmOOv9CdnHlHZGhvkcduCvZ4Mtg2RbEOLBLNzoIuVAZ0+LdgerOHGODTjay0mLcq
o8jsCWBZ2yYhHjSb7sqpDbgi/bXsYItMweED8zKO1SHE9Rn6GJ90rGJ3kc5DF/unplCGFMBgWIVz
myT6efdjS3thpjbc0UMl0ykh0eC5Lhj/jMmdbPuF3P08br9i0qKsplieEtFdhWnOnXm95e7KVVSo
uH5N3eTvwtHrRrrxTalco7qvGnJJjCYmhzccsIvy3dmxw/Z8vfDccBNtwGUcMp/helgQqXEqWUan
57A7rELBCLHvqD9ekTkFhAoouua53X/SVvgyTMiD6nFFG++ZNBJhBH/FElEtU1SSgoqsJMEgb2Sd
xGTmWMHmRLCEyD5JZqgf6bU9jqP5ux4EU85tBf6Afgut9fjDPdMwiQYoNXP5QZG17sgkf8tdWR7x
uoXnTo82hqNok8Y6oHWwTwrzc72UaJxhsBAxc6+CH4kSwv7BVXBYNEIm2nmunHLCa1vOXhMms1bf
GSc9Qvuj5LOkSaPIbj9e6XTppbh4IIawJF+b9ywjf/o1dnijfilanVr/7f/VD8X2hpp6J2cGwyhd
Q4z3c6cDxErotkPx1Wq+2WVqkOuHTjbwyqp3Xfqrh+Z+lZ8Phsq4bPNRZN4wugY4Y8UqhlbCrkZV
gqGrJ9nZFSO+nZ3f8ZcQWf408+QNiWzkDbmanSbT2Ultb0dvAtjIG9w34Wb3Fk06AKHJ6UucyA9V
29JBBh7fh9VKr2ukJ0nwXCKKiAK8IVBS0BZ5ecdaWgAlJgrfw6EKs//rgMZhYOl30GR+FGRvmZ4O
6RW4hVw1NPaOSlWmvqDOWaOXokHDBT9NQKzk51XcpfJaoEMegoTy4PuH6X26WwyqX8ndR4XP3GaD
/5IZoITWtGNfGwgZC3/r3pA3t/nIYwTwwZ6gFe0oGq9k7ijxc2o0rBQeuFY/w8QkrbGbZM/kPt+x
stE7lecFy8boSavJvWi3hPKdm0dF0ewpZsq/U+kK56HdZjuC02nDAQv372/UlqCtZesv5+/HmueM
a5RWHXO6pYyq+Gscj3HqrohdoQJVBzkau+AY3TO1vroBV2nO5DnHoRNvJdvRYPKXtDD4fZfVwOKt
J//tRXoW6j2UpVBvzCWuoBRWp3AzSYJrpb/mGEuFXwLOIT36nRYtmdte/zSNdmQIPzXFgT73NwKU
MnkkOrolU3tQ1k/yh8z4R2v1ipZu9qUKwHd/ZsYKlA/QQ8K4NXR4IYUfQGxZebFDBHIwHwBxDgRD
IXHqWfnrYvizRTbeKex0zBfeeCBfVzy/wtI4Wzae3mOVcOWPRH8zdG78gbwno2uijtPPbY5aFTNQ
S5f27x9Sv+H84T0NZzftk+iC87pmMLEHGSWwXgBIdZwwdJrdM/k1ILAZ8fjfac4j0lalgFm5FGaP
Uhv44Vk5m+8IvfSa8/AmN0hqHkxtlXUHGj2fj/cXPFu/KnlwbwkTz6HBDPMYt/tDN4Cj+Ub3iEdJ
PJYSkbfS6iT6s7FaOOm0aJAL55709wPGdnJmcqOxjSi5x7VWbi6dFa2h5uANvYGejSXCoHbsA0nj
XdzNfy4JP7RjXWVXQCOqT95jpmxNQ80zqcMWT0PxpouYuXbQkF1DWZ0dW20WIfDe0qGDpApsnhPP
sdCgjyqjbyZT2ccnzbwHOba5f5H97upiHhi2USyRpel23ENFJ1ZFZhoDI10HekD3DZGUfPXuQKyy
/qkMGM13Klp8Fjd5SnDFY91ZGTa0IG+B+JhtljUZD6SvcthRA32CXNpbNYKmFDSt7xSVdz3VWWv4
c8mqx9DxsH77ClAbj8n+TquOHHDd6t6XxoQpjyebTw0a9wKv/g2tYigCsY4sMx9XUQtjNVOZwXjO
emJI1yBlNEgR8zknJunfOT6RgcvfM8Cd4Q3nxo8K++1UxjxffW6asi4sLYfcOHQxHS9IGObgOmYR
fvPzLjLBmU68GR5aB6fIX3vBAsSbrWd3mPdIghlMBRJXdtlPcTAHEPnJ+RraB3k3gjhd2sQb2fGK
jnhSbPgZdD3z0qG6y7jFi9O3xiFCnAMLyTmlvKniJm1H55GGUSF4bmwZakdZH50PhCAJHvKPNH1D
mosDfenpsYYHa39iZa1HBOCa1yDk3erH3xwUN/6Owj1pZS/zesGPX7+tcCbVIrNYWR4II2ohtWXo
UGe21JEAxL4cBZf/8VgKsN1vitdcikU/43qcw7RR0NooeJoJl+lWq1VOo6pptjyQHVN0eXgvEalA
KoF/H7NeRQ0nIbLxZjs20H3HM6Zh77r0iMy1WkxFwNwOngjhLbTKriaw+11RX+CdcirXm7yDy2hf
6jIm+GpJolIzZYNXPbchKKlNhPHRKdgvChrtfmXOCGiKOXirdf2j9yBGMe11COIruv8rGS7TSkUT
V5ssgGhwNfbQTBiXPb8whoh6+gzFdFgCg9ze0QGX194sDUUWWYfYEjsi8xMWBzKw0Sj44tswh9xD
t/+T7UT/mqwonwsG/8eKXOIHay8gQZjcTK4fjw1O38rrBUJksjj/frZC15BaxGVcbtBU/Y7MQjXy
IyqWpmhGM/Xg70BcO16mpOhBUpCoo+iA4CMLUILA1sk9Jgg+9mvWA+iCu/f0f8kqfNy4KeWFz50X
F5d191hKT+AX/EqZBtJqSkCa3Sc0tqUS74QM+UN4U88k07Myqi/pt7fC5HgWoT6o3H/eWwGEZe13
d0R3DFxLb7CaBLVWPlDbEL0WdHtcSlHI3yAEL+03I80+YrjN4OCqsLgwCSyBji8AoaNxodgdjRtY
azty4FQiH09ZAQ7bFkbLuB3sPToUhnt+J2I+6aW/BPvsDjZkkAjqlSNsBc4KBwP6ie3H8otYUl2A
6xFojQss08X9WBcubDDl+9qvaULAD3c/7g1tCIEjqLejP9LqgGqG0Qo1Jm9Ee7eMgVwviteRKYnG
8nl3bFOEJddD1vJEkXM+3GxwcjIZSwP8/NmC8OrGz2V9N+ynZkDZXJRamS3EiOQj7DFpURkPox6D
bfZu/YjFINzkTbtlNKTHQm0iTjamKyhEzX1Z/6ah02qNMCUPH8ja0/BjcfeGExSyL3HtOZ/cXo4X
100caE9YGzC1EH9orUqoiM5vD9Mpcism8/EuMzOvJA2nLvbnQHEQRb94zjrVSryEwjnZFn38e9yU
BTT+mm2iGDj4JkTqDcPh8r17agkoVjxYB4Nv18lbEntYb44yot+7qP/ICusKeh5hVRdC+LT07nta
u3xsWaYb9/FTHQ89Mp4EZ++tgdQoWe36ISG/LedwsEviLj+5J3NqqXdzPL9xtohQ4fQtuhJcamNE
44bO9O5Q3ya/l1AWD7sWyQtpgfS3pcNqk908rnppw/FKgcRteL8/XHjC7+qWqiJaOkRsUo0oCAd4
+0n0Y8EGO/cwYtLXmjWUBvifYc2GhAqLAEQt5vpzQi2bAvjW4J1Qu37tX8JTUhRTlbEfwkJ1v+KW
Coe1XZ7jGcY+OT9LkX88NJDWcqqpL1iRSc0uzNPWR65CG5jQ11orQRwWiI7it1ixzm1O26vp+hlj
KacVLIeX9yPOQUoch/8M+v2o9ZlOsT4vmq8ng1b6/+Vz2Wc4yCFJJGvdrOgYTYMFn+J7hGKd+YsC
4+LPrHMFhWsDagQmgUqyMzAR4/6EzLdnDrnzcoPqo43cEwrnpUJpwmZGjY65Jal5VOa8j/urMCHN
howIJi4/Le3rVa5mDAR8K15B8sLQMBNzqjPF6Vz5wDZT7nVn8Z8GA9NZUszIU+e0iaIXDV85VVsc
GGYHFSs8oTinqaebfauxx0iF2kTFt+E8FLY3qpaZ5DShwIfmrlTBXOkyM+dMfNnLNIQlelURR/Mm
ndg1zWAbwPO8aw3lSHdG0R6dXZEp3FjwYsDy+iqOeFuX2mYnnvoAvA+Vxb+zx5hia56X0op94mAu
c1XCRieZsl+nGqCcrA2nx2GsFLOkVQ1fD6HAulbCmXtL8mjl4XUH7mVER3JU1u1SFAJrke2wPGLB
ct0jr4AsgGmz6dzeFcKK+FyRGUn7ru0G9ihHuUhI/ZomSmubNe54qiHg+qpcnR9/tcelsFQWDEmp
qySVuh5WYKL7T0CtYAUMDK6iXvpqndSZYftlj7fqfw8y5snz4gSSAsDMq3n9xOJBcUlzSnH6neKS
PcGR+qDMJMP/Aw0qbRXGlNKu4x3yQrVn4Ijj9AtOfQtTWY6Cd6aUO7k4oG10xE58DkTcECVdWNP6
oVzjLdXLTvtSboxYKs/kJCMSLWFUIY5wiafmBC0PB+Q5IezEERgq8xSIhG9HCsS7rffLk+UfJhy7
8BF1k2zBm1VquOdM3dxgTC+bGNFY2q9SxlrUHQzFkY7lN7DNiPQO0gME6h+WtRcERVVYAeYskYkN
mXC2e8zn1qJ2Nq7P1v6jvD5qEDbS8wE4QMJ+/GSAgJL0YgtymZD5/DpLC2cPzxjXXMojkOdO8J6n
0tFBBq1SzHA9litPl5MciFjISS5rvevX9xw+nZlvVhfQKfxtW6RTjpq5tiRoaykNEW06HiEjFd9Z
lQWjvCLh8A5JyTB0OaTPnquVMCP80BsTOkWv1ktk6kjXGtxuQvXBiF2kcx03x5AG7tn55vK+Dou7
GuY7k7rL4+N4guDRUYoZVHAI2zPgF4C5ka01IzTd2NlSeoDZGPj7yF1OJj2O7ZqVUjL9EieyXZxp
//HI1Y/cAIp5qFT0Vsq7CIK60gTE4lWmLfxZ/VxcHXSs0zFnm8Hb9dQTR7L+VDcUhVJkf2sRPISi
HLFaJwaBTEGUGb3jgiKEfssfJsS/8C523cFNFfFLJVioJ4SzbBZC6QGLRwvSrzTRwc6fa7JBi3Ip
gTtGLFvQ6xNr5ccIJFbr+Xaa1ZXYYBUklgdFNg9Crnsnf/7yzdpymhticRSYGyrA1vy7Wn4RlSQ9
6o/vIVzCYY4dLV2FjLFnE4aLFpJ/C6X3XKA4uqbGUSM3v+v+XGV48E/BFwmMILEPZP7/ryL3jACh
XPjeOBgljpuRryhrydmvvKzPcX7iGOBIrg5EhDYczd50Ykt7Uaqxf5svra4uawpyCztE/kPBJE5d
L2evGeNNjYSP1WbDP/32Cf8gQwFDm8Hb2U5dNusHhvxwXYXnZXK3mbPdH1oKknY9Cfq9fFei/fm+
tf1F7NL+83y1nHbAjfVATt9VEc2n/Pn3PkBr30LM8qOFOpoRFY9Ut4hSF+9/7fX5vdTBKx4HMhOg
MbclI4crYbOJyhGbmosVVQtL5w247OWxQkUKu5Cj84K1GXiYodN4MGy1r2GPjaFJO7w/shnymLfZ
M0Mnb+jsguho2FO89rtWd5HAOuMpbGrxrnwdiIRv4jHS1KmH3iefPr09nqGXvSbi0nef06ej0OT3
84Cix2SaGBu7XoHHsXWU3k5bFvs74Ctb9XgKvhOAy1iTbj1RGgOpnO8TD8rhM+Rr2MDh7oWx5BSb
EI3T/zu/RpLUwY4Aem8mEL7JJfUCZTCsFLWuiqN+AKEMe8A9jnFVlanQMry8MuTnKt6PLSH532zb
Ri+7kXGps/XkOY/BrQPN4p6X4XEHLyA4leJVlP5iSym2VtvXAv/j6oJFvxvyGyfvTmgzl06DpKRX
yqI0Y3hOD+DlxS1eFRGXe8Wsixu+G2qXVvfVZjqCzslZShoQNrYDi3hEIJo4061Gm2rU9ko6+C1i
BOBnu/7zNWeW4KTdTcKXPtkj0iM2rEcf09M/bb1UXH8s/ObjMD2tx+OQvYNQ24YVvja7ZSqLfQZo
JVCEU5tut0oqznJRTFydmOm9HspaH9AHooYU2jgLSf2Xe447H6tWIJJ2KfAki+qRK0+pmOeaoS54
7t6yjfp1N6eu7ORDPVziHPsX7l7RsXBqltI2V7kQuxfIhg1TKPEaWbKMFC0dNevqHgOBZU/Z0l7A
MPHGikhlQjxSUUUbqHcbIvUxYsFVy9VFdzbAZYH1cWtb5wgthYct3DCksKgqTM2mE26J5fSiMgal
GxKwJ+bcMU7Bn/ngwSfPrADt0MlJoVTzefh+ix9ENq4pwwTHehgS64DErJ8c1UoKfcErUQ086z/o
EvIAZ9RXVdyPPe8aRtlGorVwXJKskRvcIuwnF8NSs9SzdmYLAFmqBeyYwJovUcZSvPI9IVKFMh5g
p0OIwNHp8KCKIPchYKN9qrlYvBHFiU4JnfhfEDwO15QhXEK7s8zTfhxtaGAcGNUOPXxxX//74bE0
LlH3E82Xxtb7R6JnCIw09qOtkMbrV0/Y425fRZYTdaAshMytBuhqyIsLJOx64ZNggAsdEX86Dptr
LmKtxieW5SU9QnxO2zP2oGMk5WSRYnXyFRXxr6KR/kHfSEbJ49LLOas9tlpH0VPm+xAZd5jpjbiF
zothHfgGmeB+WL1M0rRoT3/vp0p+AE2gGiBWfOzp0Xiu5JecYLwcmNLs/HPTa9iGcRFy/0zxN0C+
UiqfkWTIVwkn1gRS1FKSwhFEK+JonYs7b2EAZhZk3uYDnEmvIHeZ/ZqFITlghmWXHuRQXQWwR1Kv
7xg842w9qDP+FpiirJv20zEHMjzCIFCZRO6kj14TELM2oW5cqM/YZo5ZgKTap4gtjwIXH6P0C1P8
4Bz0dptAYZoPCGXggDjZ7+xUWUVDu8pap1sAZJfLXazFYIWwtAGqMwjSxK/Pk5L+0igM+VnNwk28
xbKx5Df2TVWpbmVU0m/oOCsYuMpfOyroiwdIUQ7UeQf2AVVAod62reUv0XY/E+0xAPOPDEEoF4E2
M7/qCGq8/xxinjF1HqJr1QGi1oFeHCYd4Tmdn2PB9lcX/5FEmOGI+wcE2RfzK+duHRRpoUJpiPZQ
Zlv/wJD6/Dp51nm3z0o7n6TQPL09bgvbLgqBf46DIkAAjPH//4vwskjI6YRJKxkZ2wl2UWR80VIS
gjet3Hh8d45oSXUAYeSac0XdTosRtXl/d4lUIp6M6an81oiH/W3EK5b0eb66w2W0d64x6dSOq+uu
6No0V8GYL0/nfbgsXIWHU+gV5Qr90RTzaJ3rKfMH815vy9nY8q2yP37M2yOKlFJOvZZA+0ehiqDT
VPix3ZuQCHPdvp3/XCDtGdCVIOHOlHWFT9IAZHVhcMEMaWEaXb9p/tKouOljn2r1uyaqvJgF9JEc
NVVsUFfxWzW9ZAZXAyB8Fr31S7Nwg4JZt0Ksyshg0OF/PxEb3Th5jNXViKK7fqSYvwH2x0FRN9hD
NSBaPoJ3en4NqBa3TM6h8h1cYajJ8FHaAwtdx8pjdGZn16jmRL7e6/n0GaGQa5Y01GpDUtUiTpzP
vV9EEtuIQ0yn8NA3vD23UYd/KRAtzC7ZifveNikTHrTMSKiLfM9lXyGnWZ563E+yfT9y4rz+VKDO
oQbFaJ5DolonOIKU4y0uf0nf/gAxrSaVOhPkilZL7VriSjJw9a9179WCP3NU/K5cSiiBaAW0bynk
sLS1eahkvpLwSkoVdJvzWMiyToHa9mToaM72Kpn+8V1zRl8FUI1m7WvPNqMm4boBDLSByixCKqfj
PG8eWopVl9yqaE+9h7hKL4MLtNHgf92/e5peEpR3h/SZT8wMbnCATUJ46BlYORrVCe5kwNRgwbKG
J7md9+cij159hy4GEcYJwH31fm6AA6h8zwa/e4/aRnNZ9pvnQBcs4rCus+T2p269AEM9e/YK3wQX
rZ4tOImId1nD2sE9eCPQgS+X8xOcbbzdzobMBBTjvfcjakJ1x6g6qSNJaCp5hDtVVD9Cr/X9+92U
C7JImDxcbT+sCe0SXMuMUNmSo3aKV/tgwvD1Fg+pcYAe2FGeSCfzRgmWuhtjFaiJbQPoBrdLa1u+
i+vTAQETBGZsIi2vCpT5UrufN6ipKlmc7NMNVA3x6ZqDGYy6dGZCGXVM/Rp4MP5MZ5x8xssR7Yys
674g8k98SWLf0lBxvOwrEzyw09S3HZewGY7iozRHBHhku8m3O01qusRBeuu9lW6T1rKBcVWyBUmQ
2NbY53OviPlGprDa0XWPYZsQAC7Z2U9Ce+WcfucuSZSFPKZWG+s8dysSofhy9qNP69wHk5B/rq0i
5wMqbd2qftfJgColtaLW0v7qQ7xBi6RzLpXk4HhcKdxBHTRrgN5DquxWsLANiQFWzlGvTCS1pB9v
bvQ2ozjn794QLXT0df7+eC0R+TZgmi0+D7SbHhQsoVMRZan5BEoBrqXQL2MUq8I5MJCyMb39TbtP
/Gu6ScWviE3Glpx93gUHsJSbpgpIjlGNm/vOFykL4bquSMiUILlPe2wxd6D5zm2aokGrq64lY+jr
yXmcTlQjfmRBZWAp8UDnhtk7WKhRuyxE2NvT7T/q0JTeODTFYydM9i6Hs7fHAn1TA+tQ4PG3yY7t
mrFk517qvATZpfI6Gg8MGYBf2vSptmo5WCa2syuK7seseVqs8Vool7b4VPnvjlgDP3JfCB0s96bc
f1Ei01NeKsVVK1wJ7sBlFNaavA8SS5/HXSDdgX+EotZvUZbKyCkheHMDHD8ougLO5+pdJxB9nVau
qasDXHfyBE+SxUQOS6dVMUe9VWfosV8H2SrkZmsvZayRJG9Sk54tmNftmWIn4bRA2zYnTY1VKvRy
PlUWMXcWSJ4D9dvOkon/h0NmJc5RjtUalIoM3PwZvOk1hV3nl5M07mUkI5kGAkXiHGty66QdsD+E
8r2llPyjU+E0Iz64fR6ziv8qa4hbt+vzQEGAN+vODyWon433JgNu1K4OWbJfCPyOhYJrPJpAJ0ru
uJAhJ5l/G16hnrL4i/B/a7A8UVwcttC69mSzo3/StgXb/EoMpymRDNgQrl/ihhn6PFG3HIgvb0ja
pjVbAVXA1i2Tvq8GUp6MOVpgxDVj+GTo9WRGkrQ7IMIFXEFDyCI6XM6GqcJwf01eyKBEALogujwv
V+ygFrsAVWbPED0XQAzXq5IgB4eo7rA8JD3sJccAWQ2J0J1UNxbTcMeqgW5EMtuvIsN2152h5eKk
9nK8yL9PqRoxjjuUEclPHSnK+ZYXJJRYiGMFR8SxqILl7zfvcXkirMClPq2fQELS81dlU0KCntzs
JWd/KlBf7WnwqKfvWGKXox1NYORUYxucSog5Xv8Wjn+B7o3c9FEM5VW5W+aSm8z9y6en4jkocw53
BGxgzvPIXifiPC+5IBsTplWKcXnsPbWm7zXLwhlj4VLmCdJB+T2ytpE8pV8u3r60x3Ew4HMXMiHT
klFZU7oNqjAnQ0ybbr316k/UlL4LQqnUVkICeeOQH/LPq8KKNHTqlGUlRLOEl9u8qXJJTzkDGVGf
EO4r5DxelSA/b8AJIDq0IzDR2oGSVKLZz7s/xkENaTkPqh57LW+M1tGeBB+4KFay4NlGaof2Xqnc
VpbEOZnWDuuOzk/m8gxdk2NWlCwO9pcqmbOtaETFfJX3X+E5c+PdiNW+gMTVkwI6vmsynZQ7QbCP
yEZmFuQcAvylYHIr6S7XVfOrqZutdk1ns+goNhSWEJOgdJdlt55jzqO3iiwKyyqQg4sqpkC0+7Mj
fSgUxjhmnuAe6zPZrut3392XilAKG6attW9VMAIs4Ujt5xwC9WmwPwHX9tbN/w6ACEOgT+xzZehj
qRMFkHOna8s9UJJD2asQpEkjMuluBlGN29Ba7gIU/L7c+bbaIULvL6ZlEij5o4/HyUJ6scy6RSFT
x8CCOyAgSfckyIyhKe2jhpz4M93r92rTI1l2aGWdojyoj0U8MJOpsaAD8RYoqz9iseGixIF0Roli
DHZepuss4MbFEWVKy1yFFZYC+GJ2Hn3ObxMpfVDypKslvQhwhzDQpXkGkOeEq0IDawu9/PXD9qNU
b//2Ykq+j9uGQgwIr+e0d5HeiKtpqt7oH5xBNrW+q1FjqqqS7WaodO5wgWr/OKdEkMTkItUDPEKJ
XBMtMjkvRKIWSDYNXpQgRp/48UlcT2sNLbGRUitCEoKguktGVDXPeldRhtynwWWVd3NeBDiG81kB
uBF38u5VPKxEsgI5vf1lq5DyyDfDb5LpYgNaNo1Gt1DDjw+T+ZFq9AkVm4fBOwNSKhT1kfT9jzYI
aS9eqtOx8VmOHc06J7OK6ceOcfdXn9ny+Ww9kfW20PzGtGjj7kLPtYOL7/tur9C3Q8g+qc3FAVXN
CDZiQnWRjEI5wgus5u+uH68unOUr7WggsefCf089igEcb1AcM+UbrLbV+K7R0cbhewqCnVVcV2Ih
XbAaAqCCd1ZaGdzZw6IDQI4kNDqvdDShLNdQvO3Kq87E2/fPhUcv0fIJ0hm51Mvhc553w0Uxe89J
mUfwI23x3hI8XUWAA15JTswZizXtVx/9I0xFNRRujqAysmZwEabWYan3XMP4BaXXelM0+cF9p8cK
RnIAf3f1YmMLpxh8thXoliRWeQG1zu1W5cjGU1q5JY64X9/12KTL0zkzhGIC20cuZL884AiY3TQB
1hG9CdYuNDaIg5w46ewu3aczFwlwYPWdVBqkKL1wx4Ee77Q8J0OWj8sAAfFll6an+/NIStZlCZS4
PB+C/a3Pwp2b4K6zo/6f/4SJnkfwMo/ywwwNyW5z6Q+YeDRdeGPqyZ1K8jPXn0GoJDH9KnKoXLdu
4IBvi7DYISPl6bksqc0d5L0ugLnCY5R7TgVdmZrhGhv0+IRfP7I1v0qXvp24yoEOZomAwep9Zm/+
pqAxlpon99o6nlr4rMC3vQfSeV/fcSkxAut/Wl+WLbBGLVGxl5HlK0cKaroZLLSj/1MJo+xplKhm
RWDCCEurvCA42PWXM6lUAKkPX7B2/thmIKrC1MFwD49wksZzmPa0d8Q3frF0Kh5D1oG+CezGwdNu
xS/Y9k1OtfKtzI53CTlW7bfm5BrEmrPY3uU5X3SzacwK30NX3ngs/MRELJHUgYIjXFSNbxv2bMNT
hMXv++f9H9pgxOjr8TESdoZxP8MKInXNldGiDp6KKNZ7Al6lPLhTBcezooy+lAGidSDTBsXdOY6j
CviahXHSY0A/R0vdIjABAlDHYClDlwtKyNOZeJmuQf/frzm0p1MjYWXvn+Yi4596ZmhdTHIVdQze
om0UWtYeUJC68OyfT8E1ZlRHclTCWV0Zsg+gHJgBE9X+4NujdFcMaebNpe8SnndVfUCAX9yG6OMN
NYNhKjeJ37e7w0v3j1PIIvLAi4twFzOlIS/eoiqvzB33bYjkqoBub4sgkZo638etsF8TEMAoZZFc
44MbudQG2WLP+aZoP7FcXtUqvOzNl6cq+DOhpRM3230Uv9kLZGXD+4vXWu2xVgNa10YfGrY29Dls
67XVcd9w2xvNzl6+Pnt14fVaYzRyoPewdEii+GU/VLblR4SmO/dkvntAvsp2mqYc9cv/J86P8KRB
rkrMPNOAmFPPjLo9VMNObnaByE+m1I1Fn7D0wx4ntVrQdNaIjrt5AwPRHvvXE6zh5fsG/DlnyKnA
/rTTD/MC0wPelNVrRb34I9fgxx22JTCvCZJFne3IBiHHmKVC61vdbDxfuHC1XJDWl+HXUK+eToIK
CNflV17pNFvaGCQXT7LI7bdtUluDjH9TehQDAl9bcECU9XgeKck1ETEaWx3RPCNT6yE4BdzgWXAH
dPgmMhU+jd2iTCsxivJuv4R5D13MJrwo4x0wcfvXAp2BVIl6HKt3SvzVf4JMAgjV/VBXb+FDAhVf
/sDkuMQenstP2RBqqqzay35hABrv4nmEEV+L2VGFoj3QtV/a1GqLwOTpsaWhMDchBqMBi0jFLO9Z
xJhF8VknjhTse5ONejtpttTcnP5FAMT5O9MtTDXiGNDGddK7qrUoDIxs8AZyOK0zy//+frpKD3OQ
M9BhZ3Kl4bss6WMUtiTCV4i+xaqUAx9fPv7lYwIDl7HFKlXx1pGSTYdw0tsg/ywfQddpoD09pPjx
nXgd5BtFC375qNM3GsEy+bZd/BfbYMwlyfsjsgwVj4IU24kKS8RjLh9frI4gXVd8ZTQu9KJXuPda
G7gfVGn+kJGMrXvwhBwsyhnQXObJnEPrrIpY1XnPl+zX101zGKmt7dIUUDKIeDfSex91KhNCYbmU
RZR4UyJYqvNV4RlAfQ9LKKtSj84VeHyJ1AhAQ1KV0hz4qqjVO1OZvfpuZ6wqIIOBJutrWBVxjuHa
FKDFr0VX3G2bcyOgHSnKc6ntIAFKQGg7iDg9fqlrT3oiK9ByVB4PqeGx3y6ZelFLHGucRgE/gwOV
BLW2v1lUT//Qgl/GOD+jWPfd/C/+CfLOTxJSbQLcs7zX4+ifyaVbL7ZMZM/O1hhp9cmC2K879vFI
FpFpQJ8NyetShYzmlSEfqSooPkcQ+6PYki7Uz5e7K/Yu5GVcHuC9gFPlryLvY/Wf5pf+HINqQHVw
8bx/ks0drgYrGliU7hGmoxmsWP3H8Ok3+VYw5UZSRtlJcjR8/wQrnKGTjWazhT1P62YsJYM6aZc9
MsEuCgGqk9/dE1KzHMWYJlbrBuzaNss16p9ITHxxra5mQMwiDjkevdnvAKyHFpWCt4C5FiSOGT38
IMxaN5zvbbtvEUartNbE1NwEU+7ik9DXQBMGX6soBeHDVh9tApVeaAVno+Gk9UerJHiNvoiUn9/c
4e9ZAGTo4DTCxzikGoJR43Un+rEMF/4WDlTFNVd6mLxdg0ys9+g/bo6fsKE9R8RbcjoBDlodGK3h
rTZbgYbl5hTXinahMHQEkIUgnq0IInb45sQeUufqpitLFLLgIAlPoDj18y6StfOft1IL8Wq+Af7v
iB/1WMgdrmN7YnhawzTAo03axhlfvvC248KLRs7kxjDIyygWxeuSG5fuIUiEJqh6WTU9CnJHkOk9
TGXnk5zbMfsVHyK1YLH23zNe1P3LfZQp6S4EGS/p82k2OtueiaT+asI1rKUIdVdWzLLeD53pLThG
YoO7qxrthMTjd1O+BTj21R0X2nDoylm7T5BLJi/HyOHa6vCGCRENR1i9hbDnUYhsSwmMYgyK8crc
lcAkAB5wQthJBcS+a4xtn6LoiEvureftQblH7/k7DMzzeTW2SSMq3NxXbT5PQNXs2UBEpvxWENwX
GBn9N9jRWnKh3JwDXsH7E7BiheDqgPRh2R7seV+XnjA2Mj0AduiV2W3WiI42807bB+sh2qHJz1pW
grab2wB/AivOYeTgOK+ebceTzfjPiyq0WzhAXS07VE+79gwXZtFMMsnLK1eSB1u6/tXGOBOEVppX
S97XghLj4VzOl7GJGR9Tb9ocSzD+Wp6kYdJcq7gh0fPO0AQxbR9Pa8P37eHC98LPPo164Aul+2n4
XuSPfVq5lDEeyuP8u2tF9Sb4rdnRacQqhb4Ldz2HFM2b6RccZMGO8aKJmYitOaME6zjT4+bSw5Kx
lr17+BQp8vPUS2JSdsjOyqZJAhcpl2A4sCkN5/knCuXTzZKJzqVzKOaMRdfb+beJPz2L3ZmxsdOt
CDTFj0SFO/vo2Z1Fb1ff9jjdJfiQqQOM3/lrq/G/nZX1/fWj83vtfto3V5Sfy53jvW2MT8PGFZf6
hSpgOOEA38W/TvCDj4oqTxHoTh/ChuBoPkDiDZ3FqEvmefueL5JD4o8bqxX3g0yEm2D4RvG7fL5I
oNU6h4O32AgL+O00qLBJROmG0fe0DkzDz+G7O7cNZdHG5D/YIvdpH6h23tMs4s+7dc5WhRAKfxUS
qHT2x51KF1pQANl1MJLKdBpbltfsYQ9XWorgSttUjeHVsJXp4w8grv62ZdOQJ2UG79NSPUMyCIaI
atG4iSXjIbZ217Tmnche3JZ+v+TrLdPbmGFY2FWExBEGAxcqvBMEeY1wGYOOh7EuTE0dFUN4cmOG
04v3toBbcUll44hSTbjQIh/Qvftfdh9RpOddym7r4VbrPhfbdfBLLfiDQR5+rkLIQdral/iEzvsG
JtX5So7Sw8IK13Rzi3yRbKTlim2qiR/S+ZYFhpA079l42NmPzAAO9hIa/Kr/O28JlzOk1T1K3SY2
lNcuHhV6E6QdOYV+ZPsDaFyoYSrNUu/2ypixWB+azMI4GuoPD3e7O3iZKtvLWOgueF8zZBjA7cvA
GIYZ9DsJ0pBjGu13dXm98wLDw8hKGatR2lTryy/wpPaF1XPM4l5lIl7ggSYcIYm9Ghmi/22Craud
qMhNRgJQ7LrLxQeHV7I6IGNeb8ecObnZTViVUThjGQMFzO0/X9+Po+XlRehO0iyJHGlNCSuaJHZx
oCJsUs+30QonO1wuGsw04PElme2QieKhcD95+0lmvgHPyPvI9FZo4F/KyOe2XRr2elhaUZT9dldD
Ne7fC19uatHDsWBw9J/1oR42Gmmku+Wj49dQOOaKHOZ3w7yfpTOA7K4fMafUe9BpYO7pqaVQYcdT
pqN5D+uv6d5JA4CAEhitLVqkZsPZ5M8o7WMgGjKvLp/HMYjmzLJOu5Rp/GYDbBixKaLJzaldYcyL
mc1RuUXb22odFv8sFoXWvrzwkSg9vj2c0hzV4FZMThJUyzaDZTUJ5a2vmIuG3XI+2Udlw3tC16DD
laJwluGYyfoSrVHCGgSpgaUvVRsGrXD3tqpuB6gMAIPYJgPRq0U3lGAC0S9vCrWAWie2GpL3TvCu
55mM0lKyq6BtMnIukJ2Uti9LKpxU4ObPG+4xonx8DBhjmsdpLcUWOVQEXQTaYavjBx62eifrFlt6
Vawsp4bQt9HcXzguy6GeLIUxlBJ6QPI+oxTF4YklVDcSPT6+FfOVeAZn5GJsBaPfZbHiUpw0RegM
Ie+VGMM6dgzaeT4HP6u+rSMh53GI6QCkgGd20rxuZYyTP2/OdHTzT28blbWfi7OSdzTIJNqfvmjl
4Bl2ovCUSBpyCeLSopr+faW80+MpcS821IhHXTaOfe2g6rZ3BSSE2jpNA5vhv9vUG9sHWkgyTnad
KvYLJx3jjh5P3fuBgkypaCGCpLIS//6SH29HDxORHKkYNXgNLEu9SRwLAjMN2KIZiUSUNQcsR7Cp
jLHD/ps81f4kWUSQXJSklL+fT03aUUVqFi+3Hm/+0JDslfu79VuiNKuMh58AmCclUgaIVOz6Wv7f
HWutEEf9ZGFICPcyb8ubvZ2UW76u7DOgGKYlNNffjWUJE+Ljangw+GCPmf56qvnTx3s658uCznMw
+C01ca2RopL5dViLgXizcqgUqC60Lljyg/4V6eJUZfu2bTmK0ICxyMsCK4XwewlVFazO343pV8Oj
iFedtHSK4L5nZnKi85fMJJckxVns9XCd4pgewVE55bz6TYxhq/qimsODy2h9xFHcB0eupq/Wr0lT
IENMZddyaKGG8ccpUbVaK+FaoTc8XsrZXhLWGztAsxDX9M7Vs5170+XmCtmDb0XKYMYjIKZWWyV4
gnHtrZZ5TYvAq5wS0g2v5C1UMt1jxe5gJUWPUobrKQ6NZdMHC1KhwEf5Kkidlp5S5lucLxd8i/h7
jaFe13s33LrtK9EBmYEVtZDmY5g6cpwYsKk2tjz5g5E4B6srXPwIRFi8ixmqwXA1x8gfEkHeAqid
HuL2PO3K1cdnDVSYmxVIamzFAF+Jnl0BTzzD4HUMPBM/ZPljGUrYXUQEBmMPGtc5t7aQ85QLeet0
7Yht8kObBfF1b7zVOejA8eRuKfDzLogvj1lBOtvCcwDX5id1GcSK7bn411rNtmBTIXdjGioMfVy5
aI8pI0b3wvWsUKvWQLF73WAMQnv4Du/RBjuMm8Y2iXhbV8jFjvgQa4xwQvvPXWQaNyrgO28+siMb
R1/jzwSaun9YcAjjB+3BDpObqgrKT5vQ6gj9OtJdvI+aGRQcHuLDIixWlLbMVWtflp7eQEfG3C4Y
c5TxlyLf+jZblRJZTnARcC6DfdE8CpqlTwPPEv8AMtEax/+vdxwtxW++4RVfijPjf/3eupvRHFsF
bNPrOFQwUwmrXJ9cHm1IT4fwwm7LzWq+Zf94bP5tzPHnMl6v9znWWgDJcE5Z+skK708QXSXLoc6P
gptuy6soBu0KDKsGbnF0jFLV8UiX3mm1M/PPZ6m2qSPNYIgG+3ai02Ddc1cWH62q+DSdBDUR2maI
WnUN/x9UsVg2M4pBvbGgLbuej2DKypZTaMZEYet5DuF8VqEj9nYEBv0LwspEHZuSxB4zij83xYQ5
KykrpjlH1A7rjq6L3Ar/YcYNkUe6JzSG8T8wwE12F/6zLUVYS+vi41Ke0d1Q96gq6ocOsUAZ7q6e
DfmFUsnZW1Kj8JB+seNSpUNZNsnOs4COGr/gpbl/O/RT8fNXBd7eseF3IW0T/RJRoNQS9+0Y9SD4
Rqn/oshACDx+xrO0eTkoPU6oPwxg8DutqwljzaJeh0UdexYe8V34AmvSB8ndNm2C81LVw9GaX8IZ
aSMxv8Ein4zUcAgbdnwIzOdEpxPmIwXLrN+h0hQRXuJa0vmduFBsrkEQsWSuzaMdLdM1TcGAMmGV
uvycwPAXJVKj7jWijzfQ7k2HGkJqtk6/QZmSasUImH5tkA1h/rz/VpH13OpMKWnvxwYFbiwd21II
GVljdAdMzDA7sGhaqQ+0lNHrc7Julj75G9+v342adxTnN+gdLGfTRH+xQ18J1O2N7XoQ3hNE1qlY
8wwwwcTMdN8IgQxu152+SiHjQ+QTLoF9d+K9yUnk4agJmm1z3DC+RUxhjIv5Qx13QdS/s9eZQOFA
F+6Lq3f9brPbnX9R1IbJ1BTCHrm3lN1BRTSjD/KZ5nuOrlkGT6HWM+LPWM8RVjAxQQTEtbRLsBeK
9OWOK6ijzRlTwBNTHPBojkokkzR5StRXzbL1+OHmN4rF9OA9vY0jbuZaPpaJrfcuG8U/egL3nFxK
Ms4dHrkErYkgdLPiv3hKnqru3dPyW2RZOEd1ZX5rHdnSsyOaffNwmD+4HjOjAgWFFTkZDe3+6Tmk
7/irVcf5nskRDBl6TQvxhzbghPPA0iTTSot55AWiB0MyRlqtvcW5ISwa+28jSAYyIRmlPYxXFRBU
Uuco7Joce5ziIRV8YLobCGKWpmWELfECJv3ToGoye1rIKdrk8iB1KywYN7ZaKGaZ+Ghp3P+feXP5
X+1gKhiDnRjPp4R+pR1SDBbAoswUlXulyKeDQgYY/z+69wu7icT/nLsuQSv4/+YwXe63IDvMhmMj
KHNCTJ1pE7Uiu/6A0KPfhAwZ2gX7k1JLAzHFMuxY/l19aVVIjHlHjRg876Oy/Vt49TA+px+6Ur/J
puerv0OuMMUD5HBG4El+uy7yz0vlIi1x18WcOErxb2BVJG+XdvohpXi9b+TY+2TWe6TFAbkFCkCT
zvyJuyQm7vtcXB2RoIgZdTnYWSw2OqIMrJx1zNbCrE1CADz4mDnd5CpBGlW07eExWSRwbx0wY8z2
+Ax3u6P6RcTX8zqxnDJo5AEdX0uamhKQ6TnHhgh3ahsmcF+xOiuPhv8Khmomazr9n/S37zawFs0P
8KszwwDgfC/5VMuMZjJ4lt8zvVotLNZztsu4pwDmnCiLyg7D8Ae0TwdtuutirzBXliR9PlgC1I9x
EsQPmlqbpDSa1LsfwCNuQOgz8F7sOLEcEvVj4bKqXZzX7t7A4xa+smAufur5QJhdDOO+AgI8DZfl
jhuYgrKIzjDaIVY7KwH/TRXpokPF1MTwyNnLRmC+3AsyV9LJ58z/c1GlScDYIsbSM4cVVsYfnCA5
pIEbCKyWgciWBYwhxYhqwKd8TevFqclHVgKOp0AyZXejEuvDxuVkwLkD7NZg3/b92HzwwFZgrL4Q
hO/memzOkCwS3qT1tIWWJBfMXxlKbrmNE8TizGoSJHZ6jBWfWoxpn1Aicc8OYI00gDtiTuopXHu+
/C0Cqon3oLtAXicJ39yz26uHICwSmXt5nbWQqRDROenYEDbhiAOvj/uCWB8Gn7ExOR070rwWduoz
R7+LesZXYZN9AqUozkX5bN/nwXtVD7eQJvykRUGenJpkprQ+cMvsPlJJSTjhA8FmT/ljLs50EPFg
MxSa0RK+OKJKa1jN/kP81pOg/ZiyrUnwP/zZe4+AK4QPeSAmFvwzfeHnctpTerF3LMXEK1oXa84x
NA+GLWKyl6AzVke6q8n880wQgwYcUJctZPpgisAGNYlVLnlemPwZL3xvqlBH5tq5RCLxaOVyr1uu
/pIXkvjqu3Ird3eSaktRT86n820UYaI9V2B5QkbBeW8PkmOMipAz+RajjSNvV4G1E7ibg0gBu1bk
th1kGqmq4/azeg4PmQHS7AKgrIM4to/cwQAKxFM/YwHaPAFphnp/QnnJv0ULmlR3Me9PLg/Szp38
hRlTZWYVjr6CcDMdshCr0Us2erqwPwO2FR6KUudo4g4b3JRU1kECyhQlAYEKVDc1VgIMmwT2YrbN
tlBjIWzgmdiOywMAF2GTii/PNohDdUIvaEi1jTjSufcMqHPFn+EkCwdaYVOlBNk1/OcCJsswsH3j
c1Fk8JSqMKYcAZAU5EF74giZPomvtzOg4e2jTYSnab7fRmjYq11XnfpTpg2BwFOvzzEr3/DtFrU1
YIkjhyFok/hvWDf7B0TW/E+2viwteYgvJPZLW59tpeyfkPMvnGavQCmjHvmno8zX4bikxRKQ8GNU
PhQTo85kIdOT6zzm9IbG3eCZ4L8lsABl6wad3b0BdMtdSpCWlYjsWTHNgoAEWJaCiPpMYl9GaX9E
Bs1li1GuO4QVQDXhuYwTEsN1NwnHVeqJT7r3ZEt3P6AFSejK5uGlXM/yGb35t4XNIUb1Q6WivVUw
HgmKleRKptqaXQ/k8rjQ9TS6LOVuvlxFCcW1cZMRBfiAZnoWBPFBSLAq6STIEwiAVIFIZIxwgffY
7roOszMJmKUFQMn55yB/nTMEmBrq/lUWi2L4Jt5ivq487W26oLYhdhOI3mztv4CoNImGFu2+D5P7
HDqRi27n/tQqEg1BMaX5P8LGs8bK9zGlXQZZFUYwzvpg8wAh4nkHbdima3ZGLNdSDpJdTAhkwZuU
WzYy0tAErtklYpTzN51JXG1DXarnOFPj8yYzOq46dqu6LtSuj7+bz8cM2ngY9MSajQWxiLQd6svb
gMBmBlmEySdNiA3N2hvaEHfDpUg4viuim8TcIi+3QsqKIe6EW6Kj7eQeAL6KeHhIHEthk295X18W
pETYjat3dU1TzDv9jqKzenOUZA25S/oq071Dp/uYP2zcm95eE9eU/GaDYjoQOD4TXgUUVxnyJXFS
dhuar05qxH0aWfRjIxqba+xlndmXtDc0/DY62ST0zbNRYRfMPaih6/pbJzCyytnuAFM3Iom6T3TB
Y7AqZN7VzLJ9tAndcnU4bU1a9c1ymarQzSHfya6cawl1+9YWkSpcgY0KHnJqyUgFOVILLvtfw2G8
BT2btwdRSFbYmKu5r4rDVrCGqFN6uewaf0jpkpgBnQlf6ezNklm2s9PUEEBFgohPQJV3vH8x/Xp2
1FuI+0zdV38ZNsJ3LZpOJsDnQeMtue8JsxwPZjNqY4KcZnrLE+XDsEsV2paOXKLsGYatbndSQozQ
mlRiF3b2HrC10KfAPChcxloi5c0PzJ6bjy4wW8ueBwuRvidnkulsrkI3D5sVx3spyfk3GQRqF8LZ
srWAgBY6pWrZmOEHjqTLdwxstGpkatFoek8EZLkPI9HfNi6FuC2a9SAIc4/nEzpIBO17bXc4s8Va
V2NxceDQD0I/QXsfhZmouhZofY7KE9R3Hv/nle7y6ZG31FNgdhOFKBFJKaGhDgrlKLvy0GQKwXdZ
98De4nI/5JYUaLTtNci+0yvnI4VcpvtwdhPy3ug0SoOK3VIdf/Vg+VqJ99VoZaorMuxRdL4AKY2P
yv488EGJMT0El8o0thG/rCYTLQ0gy49IsAGMkGwjYOU/IgT9ANEHlRhTt2EWO7ZLE0dlonwMTgha
viugkeU4CqFlja9kmRGKCVU9hgr7Qgjqw6/hK3+6icKglj09nnupz6vLjAkXWxBmQQGTemgC1KHo
elL6Mh3gadBj2aHbVAn1ilA2SiL2DRv94TCRrMzIEXbtW16EwxqO5u0xdgiFITjs88UzBiA89O/q
D89XyifrhIVxFwvHKBCDdebdJGUfig6qkgiQjDz1ZLN3wiP4N52rrUBCSYEpiNbKZB4P8d1MJCUJ
rVqWgVSUMN+oJuFtp9y/8+AtfxWg9uAvTupcVJCik3hTMPFquqmU3nPJiOGjwvLXjwBEAYjU0RM/
1pu/I5tGk/SxLBcdS7pG77p3f8yJtiv+AG0P/o7G3sMMkWl5qJwmrycdWMGlUFjILskT/qSa5O+x
1SElaxRxlSTi5zv/ul2Szr8XHedO1k3sM2WzYyhWQhsvSjTyoX/rltzXDncUsQG6UA+D2ayYrRGC
g1HzHrSqycj93ESqshIhw3rsXtf685KvJexQmUvS8oGySY0F8Z9YSM9gFqrPWVvPHdqhHgshiJPQ
GriWTy/BxZIilXEMnilIL/dplPOBwGQ0cB6WZhl1ej2cZIW2czHZ9UI45LaeHHBXxu2fmfhw+URH
5tYKrRHdPX4aiOUn3J6O8VKHISJw4kRE8nae4Fh52FJFpFpYUX1iLIs9uYl6bHA48wzJI56UucOA
DSyeQztkSGTDMbdOnCaROMGVEx2L3ujpTPyL38zBgc4ADoChW6QUDHhyKAqd4bkkAnZoJzdj0Zjl
JJgjZaZN/3F+eP7nmacUPaQoaCoUeTsdptLj9xv1a1IU+LYqqtk5deVC/TlFaWSLOqHEo87QS/AN
QxndvxqKNbioXt3Df+iRuM0Xzi1SGcsuxxARje9FHcqPK/NSR4AYAl1/VC69XIXe4+Pow3ifRup/
ML4yXhvSBpOjL1lRjfRNvBmyTVz4Xyd/9/mAxoKxWm0y7q1Moo7V0riZTtA+rO9yII5kQ+TxspgT
1Rt+0ll/8ryD6i1LlhrwOsKJ1krdKeZVTeYXuph+MCJv+vv9RoTR7L0FifLCyYtfdZgrX18OFj8c
4ev5uDxGVkhV8L8LG7TutHXBxQVjdXv2owes23PivqroDs+bIf++1T9ZOlLewdHFX/QzmdAR6SO0
TGzJkv7ECfh+gVUXli+gpCuXyxmSPTwI5A/VQpxWCORvU7tLW71Wba8EhVSGa3IjWwD+6FZ77NPe
tQ94XF295CgvXCleAM0LL3FrYoH1IFNu/McMJlR1mv8hJLVlC/dgYHL7kxrP0UdI21D05xMbQWnt
biUwv3azWuFL33+zETcAcsJPUTAhty3j6qxji6c2wVWklf/aY3ad67tJ/FjQA4X9S1OUkVAjfrI1
okj5geMrpCvV6GqMv2heHKuaoHxTgup9b4VoRb/mcBaaWmPf6v1+w8RD1JcLA/4rYDNA+njnaCzp
wRoLk4SqqPEb2Uqt+ln4LL7ihJRcFrHAaHu6MV38dccP7EYfVOO0ySMwd2CcrYvVpSAhq+70OBbM
MMAkCIDe2lcClWNVjpSZ/tBLy/touJDC7suuVA0ed9xpfdnnTPl/72uxIQNSdpnAMLTlwjnOdjmF
zh/kCeJZyXa734a6K7t9on68llQO65eFZoKPjG9fwATb1Fmgft9gtQRHfU6oDTLwNlI0sTVgfEzG
M8t7x+IH+x2BFm5y0WX0xlEtr5zxyWNxuGRZB4Lbk43o3reFYteI0vFkFjw87BMKCQPXCe6Gh1Ip
M1Id/YUch2uf9WfH5ic+EjSqER6LFGE5P9RTaebT+3oXsOFuXRhZMqSih5Eqaorq1g4AA6h6xHeC
5va1OBG4JcFDafjqipgsM3xAaKV5BUbQfjE4Tl5tatfDPqUPwd4oksSKoSM3oYEMoLYajybirEky
yO/cq79p2RijU+Ucoxhdri73pbs+TI/unv69jmshV/5f8f8hQCdD9XtWy+cwSu56XpSHlOUxydIs
W5eLrBHjvJYV+47Cg6HCLjMLbb+fCcCQNUu71QmDaYFP0JkdvZbneCQ+PYD3fFzw9lCcR6EavKh0
Fdcacr6/Vm/cxqOCvH6E8OxV8nfgwjIOc9sYKnbSB//CdAsFGLV4qJ4dZ3QXsP2NtoRFtaHb/qwd
AGWVXdkmu9cJsDK4ODC+5N1Dv9YVqXHGMMMs0T2WaY2fvKyV5FuU1695A9C46swr7fE95IzYnODO
pM2IXS0El2d6H1EuP0MIGs0aFOHgM6F80+4+TY2as6+ZBsUzl/E7xc9yjumxIIiSh4losyqNOfD5
QUirFVAXUFJBqo7xvffUXW6rnHESWBeAv+E8a9hRb4O2AmCxG7oFuN083G17AIZ0bVeMYVMbKpxn
6FhoD6UlOyBCpkSMno2+O3uxt8wlKpNdmyh6KaiF8OdRlvjUY8HqxhWocRHyg6ayZLSqRjLMCAFZ
+aI8rIn1YGiR8mc3cg+YpED5pgeIyNjWMrzbAt23N4RfWLPbOkIcrRkKJ3a7T7+Vh1WGO9w8rqWj
+v86EvJbQRCAslbkEM8n4UQlKy9OmWneWp4MHn7PZVjvMWcG4m9VeCcM3rhDC4hELMOV90dWlWmx
PgjKk4ORwpsMUJLgbCU0g1bPfs6uWheiQWNHBXEGp9V9Uz4XfGuiihzwUha9C+x4OriNK6s6rVFp
/c44o2hd28iarSLvUdYuEJFpLRS0/N6585uacCMQscTbekI7zpiGG0R1JSoiJQpvakkgCma3tFXD
1B0TfB6z3WCIMfQrAwzsis7siAeEJaiIK4bNJon0MOp5lP5EEILExQ9jqkn8qUHmToILssaxSEtW
4IoW+Mh+EmWPR/93m7Gy1knQin15Q/1Z5WoQm1bRX72dGfTl4J1zdcUwacQzFqD5hbndqAV2zt+6
/bsUSiBlmcVAraY8xwQFpsPGx5icy1+x3bJdeRAvtHT1j9afQmgBY+OyDNNbSKm4t9Fcr++kcHuF
mFl9DeiN42/+bGg5ebaEg+0ZJu5sA4HaU6AP5gqCwZfy8pfySosNvB5OmfxF4lyIy81MCg/czJOq
ZEj7DRawufiHTpqXMzKPOQERHHK10z5GcLgJUgPcUYh4gaXB4i7OkuNkZ9p5JS12xtbnNfc4yMEN
J4ffQXNm8F+OyeVmI8rD3orTK0+M6PwgYV3rZsGTk4mTByOODjJt7PtyEqOTcSze1A0c3m9sK+5v
Ux/1Dg6uuBcY/pNGpPP1yRR35C1H6fzPH+E09wfe4qlNfHjHd1Le8W0NpUN5+kDjjFUZcTvoldEt
naQNWmoTbym9Gh444ftN2Rj+9qXDei2TNtONOE7kr/MrQdjzoouRmLch7+uafENXOj/GF8B/ngqY
qp61nnek6s9roDSheCa5gTsSC7Qo2wpKFZAA/Gme6TVeroQyhGptrJ1p0kK0y3JrTmIH6rvkFGMN
7qscGY83z1NAAhgObA4NttJ5ZAV9MukU+1k/xw+jNHSDwK/dGzZJd0puj20WJYWC7CNsw6S7LaGS
GUL9XipxN6JPu2IrSwXFAoYiHV6ZiA1lBKss5Xkd8/hlUFWnOXW0X203MDJPmGaMFV0frRwjcxLz
iZS9Ap9QG5hQe1uIrM3USatWWeGLxXoqTbqFZJwoFOfM88bBDM7IKUYslUnpYzB5UJ7jNh1jBv/q
jVYWVyRH7JLHh+ZWGHViy19c2BwnNgk1hk0lKpgWV4LUgCLGlvt6mAz6huvIxiYN8P0Se2ctn/lH
dSGpKuR6KpmFNqCSx+5XNNFZlMbqVzPETL8M6vh2uJu8Zo1KPxouiwFy45D/IN1C078KBeRjFoa0
QQtocKBghKe4r5Gx9C2oPO6HY1MCVuUR0ZrpGN4TeyuYH5YkOBzOBkBsSJFOqf6N4tyJIfNCBK2M
R6e+NIATIRRmm2URG8U/mY5uegI3ucWhB4MkqfKipyNNZ8uPY87BcRwt7hTCxo6zQ2YTWIsvVSAc
GBDy2ZxM6qguZL1UYxN3dRu+3J7mHJoDMevV2MeckZsm4fh1RiD7f5vYtL0xp1n3wCeuTf1ncYE8
2lWMs9YpMIZHEJnDrnjnpouxnY6YaVjEBtzxFx5G1hIKZXn6eKNbQpr9X0KpYQpEyrjcFkt1mkMB
mBnFGEnirVU77QPTP3Z7Nc29AulIShZb4wJ+uLp+dJFco2QOMpRKc6wGYbfcFB/IyWMuj5Gay41S
j67W2ehCywB7MAplyHhhNgDEZlId1hROrzngtzm6D1nVTXrA6zhmBez/T/NsL9k5XD3BLqKdT1Y6
ZuCty58Jwfm1nb0Lb2lxW3OGC4n9i8RM2ALI00gu5k8XkGZba6OI8qtIpKx4mRedfm8jAn9mEbba
sqrrXlHUyq6VysEaxbD71us5OH862RaCjWHE7L/g/aPijS+XW5UiouVkMGq69RJzoksalwpvdtDC
CwZqjzEOVjc8wzSNvcqORfVvH4Q2wQnYoDTPp/+5CuJk2hRcg8P0X9rP4/loc6K5cU00Ht5mrd4e
IPejd1IKknq2ld6sXCj+I8+x9n9uGX6vEmSSW59qO36MeYgcWNpa01dFNeO6Q8JkkCiKo1r9U6kA
4herx/Sh2MMnJNPwMXI1IIH/erkPw6FtZCVvwZDIDyASHGbhKKCSIx2pwZmMxca3GUQ5DPSnLsMr
1n95sB+B6AY2fH3iucW03p54q2uHJgax9JCFrv3fEO1txve45QBMUOHuna4lAEaCk7tGijYsA9VJ
0xKaL8tqivj6NjuQxFWeyOm37nhEANJZZYTjBwyvXkmhvCfvYlUtSWvTlSsVuYAu3zlWgPHcyDRX
gNCUUfSeQ0eyGvdiyu8l7cYuRVjsQZPC6C6qjGGRrMl6Fh6RlBANgfFqdoCB4DudPlq9RizCMt22
bv+ZlfN8vmiOU3iK2jSJs5aIXzd7xAj6xmk9P6Q6AG465l2L1f0eyR+EakzdmosA6RIfSf/7U+YH
CjYFBJQSnM+ZD/+0lH6F3vDVlvkR3HY56RG78/JvAnRXjVd3gwTPbgFqYFvII3RK0re1RBg/IqIE
IJ1rOfk/s+tgUW83vyuEWPyjwWmP4KNpVpKYge1lZBSVYUEUagKVYFIE+Trfy3xzm8KPQp1pz5RJ
zpGZuGJHSBMNp6S9MXlvWO98/X/qsVCkVL+s06qFg2oDbE25e5SIPBzC5lJh/c0tpyoGtH4AI1el
zF6ISqDC9+igjJVoFG0WHxg4Qbfa7y+EJe89E6tmbN1gnX4Oaigz0Blb5o3iZs0q1cZ5tYaPenEh
BFiI74FELpgShIY8b6UJTfLRFsHsUJdUSYknsHvjaCbUelG++fgY1YFBEdJ//iyUjyq0xj+jgTtx
GvjN+A9Dmglvn6qu8sYy8HyQt/FYIuGg35Tp2pzT9UP1hh1aW+TGccYjtOYAbQLyT4l3GJv9eHd4
BnCalDs7w8MVERMVES+biqmjSEt5mTjjaTKNYZfNuFb95leAE6yOumptEKAu4yS5d3ErZwHE872f
RMh8i0jOgyJUv5fV8cz54OJxjx4511IzJorW8tPgB4fHiWERWnQ4f69c1/eAS+dU17uI2O9kYKgs
1TbqqMJnN7oMXD4ji4ubIeUG31/bQH4DF9qZENOjC1S0zNedjKQ1UXaEnuJPWuoHwGSFS+KK+5Fm
COcBB/23mlfbLtX5FbAAv4Kh2s8UvJM+sOowFEl+jDsgV0uBjPA5t7nUMl5Jkhb8HkgH9TNzoagi
d6LxRVIf9Jtrex08JNCTNaLJY0WGCOUQ5X9nFI4uZTUfzr4nwQhA5ssr3hzwC/h20m1VprYQfdmm
2TMk+iIVT11eClUdtYE2Mrm/smLkfyXARsqkX7jdJ3/V9bY8uXjblS9cWKeu/OV4jvuj3FgPbckW
IwF9LEatLwqDfhOcsh0GzoqYTjTh9BrZ2ki9xcsQtfapby1yXu/sFciLYbmr5w3hqoY5tM1BEjhX
digZMsosQlNfg5N1lssts6hxE7aGSueyrTg9gxliMiTmAb2OFGZzdNF815cIAz2uxPy66RMMdYHF
Xblz0njiBgU9QLmlspkzgyfyxUwUb6w053YVEK6V2pFQ9A/3ieTxdp396LAMpEzjoRgBycr4ib5o
Y4/fN0An+hMlaRMp3gVm5m3QdAp19wXnk8ounfqLx5HP5P7BFP+XLHMdsoEq44JMdvlFDiWblX/Q
MNgcdW3zthzyx81jE/+3HJakFUbOJc8jzEzoo+OIavVxuWmzO7qBdeVbjxVp2P/epztW+ldfqzOI
IsBtaSOkUf3byh0KbwIxqvSVREc5KDYkDbXHl+7WnJVUs0BIW97WZPp32OXp2pq9UzIZzzM2rJJc
/+IMjUDU0zggfFNUUD45nkuWPMehlDrm88BaoFpv2JgpPhe91SKuW6gEvE8+d0Tb/7XfXL5omjjM
BJE4geMamL93JV6c0pkMPyliMa4uSOFara5ePxnsSaodoKbxSsvtdB4/noshMhJ0PTbUBWbgOtgM
kniA99FFwMblQH2ND4lHfRz+8BMfA6u0YI7UffJ6Ud2j/Gnw8B5QLLHS/rGoLAI5/B2YVsgA+myD
Y43XqGO4W0VVAkOEdpUWbwTcIJ8qIKzRpWUt+hBNrNtpfjgQUVAKy0IcztAqoo2CO49KmIKQo81v
Visi3IaaM2Nf9kGOwsZMczar9BmlnbTopP/uSkrmnp5tdTNQCotIFpL+8zMDqwk7U3NuFdUy7/yL
mR08wBVwheE47r1fxEmYLyDZSoE+rzAs/p04AvBlhHpvGS9TEGsIGryyTIG6OSqCbNdUwpOCSWV+
NrLepRUmk96UFqjA98/k8n+WI+68yaAwGefCtpQZJJfIYEKz79cuXfBkAgJ1rPdIJf/h+ED9H6do
ZHipJ9pquHCzxPBbzKTYY51LlTQWYQvPpLRUouVs0UnIr+WIjV7XJhFEPZ2KOrkb8e0Gu53SB+kd
kzOJuNUbwDkawZ78f0ckmaw9DJNok3jRwD6AMhzl/0z9i7dgdNqfhXJDyScSoS4bNRh6I4LAeKrS
+IXs/loydLgv8SyijRMpv58q1IBDQ0vL4m7ukqZ1bI+XCMzVlP0zRWB35dS5ADASJIg1E+cA78QP
Sac7uxnNcxWsox9B+ksyy1eJbPmXU7Qx27pYtNA94tcpnj5UbrmqeHO0Y+twuk+Eu4D7S/bLjGgW
S/Id64LyICx4xlzxx8GZ8u/zCAkGmxM+8p/P/JCP/fj6zYuTB4f2hN5f8P2RR62HBo3UC1wNf+rd
BbXHqwm9uloUvvsT8BBz9XumiaCVAe0DY/1jiGvmHQRjQqEjyZyMWjPAUM0PiCMI4tB+DnMcxFJ8
+PtmfmT8fYi/VwP1IqnLolsawcysGLiJFuA6YCeE4Znc5kaPWKG1FJZQhzee26NCRwA/M/dbdkxo
DUVkOYYRsRPc7Jrhhk1eJozKl+0/ruPo3zLzbx/7X3t2OPm3+YExqyB4Qvm2stfjK/qZMiufujgq
BbWAbPsqQg68jOt4cYKM1bCz2aClE4N++zJ0bVbpu8D6Blct82hWPJw5HZTRVSio55t8nFMmqnBW
4W4d49CRc5m8b1yMcaxFksibTazzEWHtS6GpAAax+VE2fl1mrHkM1IJsK1SSl7MKj/XTQ/KNdN1C
fpcZUChK00w4F9BKVMo4Pz04T7K5FZZ5ucGHV5tSCapMfQQ1lzhq5USEFVSg5GN6lCzNRGe57XTM
bGOlsJGCDSn59kq+GnNj5jOarbB5qJ5nF41j6aIVPJokXqN1gZTHBX28wJqSxVupixKYXk0AnlNw
jqZG6quofWl+7IV3z2JwS96hLKLNMK7QS6iZpiGwFgPe92ViqV5gAVKGHfDxS2xXyOdDjDQQZH0W
1gC9Y3pZWTcIMd9uxxtJrzUmYpMGMbMhmtE8Ji4zl3y4lZW3qdfQqCskWKGtHFyNBZ43GvMEi9pu
S9AmLJjLPeHvq4Gkn103xNxWDBM53ZyY4vZQ1vimOZ3NrCYK6mX9NXPupbI4GIHqvvfEMOfzOzqB
oGPf/wtATImUsrUYRu96mHDXIqMh+WmSi3+fu8okIYblD76OBsB28Kd2Q4Txsi466phyKo6sTXXZ
ccMmJLeo5fI8HzKg38UGaI4WjDiXeBVHosyja+x0w9sgCWvzlswrK2tHTGeDZqzaNAvqDUJ3Otfn
7YKgdal1Ch86KPvzNgPYAZ9Q9HpouoxbkvnJME4+X3M00OzTsOnTX1kZJ+4f9lFO2hjlIGk9xHxo
CiiX1Hqo04DOBIIwvW5deqIwn7UOkpYYKtWZqyUbvjvcsdyJ7eDgTTPdPlFSxn/NGdbiWrvSUvJ0
WrVDnmQy+QW6RuMZbavLkUEBZWweK9RTgsEKKREfiVhODOuPWdsooc1BAZqrObS095iQBVShLS4y
futToXA8XtfH4REYO8qgZw3qNjPejAjASHgKVxXP6cNIpj+b7gl+2bHl1BLC8dmCc3TCmqKHH6Hv
/giZzUZ3bkNR48rSuid0WsbLV0T9LJBqbvDTEqPXvGx5q6xmxZAxiGlr9UppWSsgeU3u0VmElnPp
v8KTwHPtfRRB5cLrS/6Lc/8YJjDf9TNj7FejNj8jIOiS7fMGq4orDS7SvT7/dLG9rbZVE38pGanh
JaTLxvN2FETQFAqhiICxSb9l+xLf15SurTniO2qSyjNCJrKq7gDU06J+vZWAHIOragHy2SA6CPn4
fkU+qVEaati5GNztsO6NCscze+pWoRxjGaw9zEcFhSRRFadf97AqcIALUbwY4xstw7QB1T8wAp88
mK3Fhlo00WTmXmwQhjr1rJ1wF9n01kAEaK62BGRgk9NCfw4jGLc4Wl2JcjfMC6lC3LP3Wv+kqVny
1a9GX9n9eLQIb4+u8FfBFlxBU0g19MfZi1TGrk5C+WPaDDSHnQFyYNriFXeKRQc3stPxD9gU+Bjk
AIIt3jxpLWZTkAmDnG5XicmXb2zRX9fCh8/SVAM028+v14DR8xXOb/JAK/oA5BODqdfaCBWU9PLd
rf7hdF4PhDIPfVe5mZJJd4KIIDIRFUwLak5skyPBGN9QqnTP8tJo+Vkci7++LDAJ9XUh6E+K+rMk
RyvqU6YJ72dl2ex9vwwXwgmW0QlCU5a8mANUL7lWWffuGberDPxWr2WreejvsSa/Edcq4d981pbd
e/rvzzQ08plUhGl6MI36rHqolBnkP5K3BR7NYWqVV57dijPHiF5h7+jWlnMMn7tDpM5JNBnha3w8
Gh25X38PVUcEfCm9IlzkPMwjmXXurplbt1pa68aFiVB/YdXYlkCYgkV04jemfGpyqvxW/IaGazQg
2s40qmFZrLdEerVbiLWJFpd0zBBT6+kAY02Spqjsf5X3ZwahZjpFMJYzn/qWrVYaXTChrRUoOs4a
0PD3uHypG56yoWNnepAwNTMt4sw57716KgAQquO2ToZtBJ3BAGuNP9T+tV+RO/az36nj2FW2ghkn
/VnXwiK5XUn68Sm+nLIx7N7IxvTcXn7LK7NlvsjNAjPv+27EZsQz9aG0Ym5T1WsiCrtlt/s06XYg
/GOTcjRV3HkoC14CFy02BCtHJkEcyh95zg2HfZzlDdQ4toS4AYnuyflu0/Wou8W93oFou6PsaxpR
G4NKbjKrtBD1fTabEAdOwoEFhXkVojiUyyHn+Qtlfm4IIodYbYmAvgckYxOiQrRJB9hpDtvDgEaQ
7T+oHqOgbnMxyTyZnRlamMGWu50aPZz8PAAWfq0LilN7aSlaBYKRdCTDzJUHBJ4ei2Cp9a4HPl/n
2xwCQvk2G/dEz+xqQaDMFftio13GsMRx1l/DnxQ1Alq2crKIPG3ldl6Zy880cqHcuwfQP0P2OJQM
uAm1ku1VP12Zd0NjSHObj3F5VRCVONfU8HkdePi9YSR7tG0VUuBU3bGzUE9cVkLclQhL59toWTAG
YdCywNEA2KFhEm76fcYAZ1J55zNtvOvjJTK9Qu40WJSHOe1GLAYG1/3QpopnMbFr3Y5YGPPoukU9
0JAs2snZoeMYfQ68Jt6aT5RplGoT4zJ6fhQgebAvmkyLBnXrcx6rktrsbxzLw58HVyAlUeYmnbab
5OdOqg2a2mXOPtkDp8wQ6uHiS4EmJHKTM0Iw3YkQVcN+2U1ft47qdDGu7MLhboT5gZxAfZNaXGEO
vDBlVGLOo4bTH+yL0GP9wRI/Pv2PzpJ1dFYAygNTBS/1wcrjHIjprgzzYbKKt69G23WKks33P16G
pqpgvXcujLEqahkW7Q6Q7BD2N5yJmlHR7wd4aBIMh1GHfri2/2u+pIBlZUw+uNIxmpw//ni58651
gcEsYUTJhMyT20S+PwTdGrKTawv51XUFZohtfPdLNOiCesnDl8q+qzTMFtxRKMC36hPAQDrafO+R
kdsFJytu1wMPayNJasixzz+TIX1b0fylYboRGlUorYNceNoqCDMXHDd6DZCfSM1850esKtuzxKnp
X75hgbwuL8MpCD3bSR9D3b3qPgN659Qbq1xh7gKF543BMv9Gjv409QGROWjTUxRnlh1QDt7yZuv2
vDjhAk/5CgS9GvJjMJ/gPU7wMIf89/j2PX717evti5yM0KlGdssbJDKBbYocinwX4Isxh5dj7/5E
RfkQCfyNCcG4gX8YPkgfksdhpqNibA4AtMWd153s/Zyppqc/zKYTEtYfeuuaBQldiiuwbQqLvbQy
W6Z9SvClcEW31uBGCvT3shFCI1ZY3F3RKpjZjC3L4t3jy7TDWRjXZQo7UOY5Bd3D8Wdh0WKBrxxl
aWJAYLu0AeGqTzdTmkwvxFxoMFe5zixUaT531mh+Gl/S13vuHhbln0MSpYk7v/c57vEIPDUPxDm5
+MeTKA0x61ncSaci6YdkQMwOQQiCWaEDtjdmsHnZDV2UVzhCoYP4qZ/TUWxYOwpkxAiOHae34Mn3
bYIZyAXkipHsbwOVSQtOjfkIL5u0MGl9cgjNC4GThxbtRSbFiv9PBMtCdJUbtC45akxf+F7vD6Tj
AvGk0892x+ALxj1bGEsNw86AJOMmpg9W+gS39mN7w4VWSy1ml5Gjd6iwSHl4Nfh8HWG8LbtPbmf4
YsiyN83EaC/ciDxeWYvJx5lzBD+z5g2b4yaSIyux7UlsQA5FUfkJJfoE7HK45vfP+maWzrQKBvJe
7VZDDNYiL2+m/C/MMPgtAmBZC1lO/MxdAilp++WzgQkeeLPji13ZkFbekrL/YneLBlFk/8aqC7bP
xzlJd03eveRvyU+64+Vxi3VZmg2QIpJj80E4IQPGyIHPSzdZRrYzb8qpdXeidC9zENZFivnNeT+j
4exlmjnW+MrxiKktQTq2NsVykRpDAQQX+Wbc1T/McgIfDMDJ4xOLpbTVrAbBmwPfaqwMyKTfBzRh
XWFYIuJVBB569p9jFlfX6WbTASYCOKVmFhXD2jjr03RKQ/R+W/eVw3+1ch3+ggyxGgXYEWl3syud
hixKgTvmAz10U1Mc/hTa8kl5LHOdn1QQUob5bYwCa7ND76LZe0Mive9QFUFrPZ7wOgHOjr4dF5ov
4/9n8/PU4ca2hM4rBwiSL9ca/OPPX5LJrdjK+Y+o9xzbwJLYcYhURTbsbGdDWFhq+Ek0ZbBN40Op
zumiEh5fxOtV9nD6EC7AM3ON8qZvEcPGMS96Rmf2i/i2yTZ8BA0+Di6m8mst1LR7ghq3XV7YlaP+
NzLRE8sJzOVzPObDhiZJz7jHVMwPYOs3AamAMaWscCJL+jQ9agNxVVnRNCvvxxkOEc+UWnZcFZ45
MJg/RO0gakyTxzqWnC8YL1vL/XqYViZuxGcZIcvwOWMhCmPGApRul667NX8KimmNZy0+jsQdxpfU
ZLzYJJjYshsJ19rQCX/WL9UYPkSxrNV8XMrxubGE0GOXyUZ2IYQCK3Ni7ublzUuL75U3P3yRQSut
Iz0OnG0gondkl6cRA2Rsy7TFZLlNL3xMYUxxitJHRwo6q+NIfCA43NKvK50WgxqmXWwpTXZgPVxb
Xl73z7Rct0TCZH52s49WIUmchdQy1fslZpld0c9nixiXriFsxyerWuRlApmeCTR/mGXLFH8yDs/k
4LK7Gc9qrp0/7ySNLOsamQL56LY62Ss+HqunnWfeTZQuEvGmOojA/5GWorKScxcWdQJE99/kPt3z
b35IlQwyNKBDhcE9S1PYfL+Qme2Y5f0SwP5Pd26K38A9qT7ZdLfBsbjZWepa1F1h1LEioqZdoXc9
ethPcazGjhvIojQ/SL0SkjACwd474YkxyumyEkSfCX9XDLLKVo5pEHR28ZgUqYtPZD54sKHcM4kU
mHTOJYS4lOPSbO4nCHYpHMnD5sipTIyhfojdAhVWh6qDKNafeRbb7vj6VIjFW67kSkV2Tpu43Xcr
yGkHfHzSFyY+p2fYBfyOoD2mNoz6gynLLbbbogqQhno9GwY5MhTAGPgoOYLfW83P3bwQqGDbOTzr
7qtc5O4Vwr+FUpD+X9PzgufYnX9jUfT4vKfeh5C68B1wDkHJxL5G6/Jsf8xhXwAV64zw9YvCe5hF
gcDWevTejWmNUKiAYVzoq3iweT+HnRk1do+n3uU/NGjBwpvLe09DozOckM730p3ykplGi5SotM4N
z39B1C6ddllTGMW7QIw/OvXaVDpuWYSa/goMF+OyTlPFsQtUD0pBrLf6dKE96fP/VwNdhFodjcb8
m097W1OqEN4f71CR9B4ur5D+8iKYDKGak7D8PyEhgTJG/G/WKdtabukftICWVm0VmDl5zNiCxAjm
Ug1fRolBzcvdwm/V/J3o30Q6jLz7WfgoSbkGRSntLqnFlRaFFC6ZS5YuTRUTnrZmmkVisvHkDUSm
pC50rUoiS5jGRlzkqQuwAmThECUz+W8/3PAgWiMWKqcSO1YZ5hwAqGxPpKBqFMLnQSrvL+1onzWF
rXz/ysixM6g52PgSbpBMYDlWQ5Q+hH+jAoucEaScllhBzX59UntcPjDpzf6VHZM8AZdpU4jSGK1G
j3TT1uxfmpbNeg+ZQYhVhNkFuzleO+vC6KWD4QgmUlHaBbBV58l15N064cInTGbXT/j4vfzzX4G+
L/p7F4AqPw95JmLYQyt3kcnZSsY1d9x91qEdm2EgNUWtfEqcFqZhsDIfmgkqGIDXq/1wFeC5mgSp
bJF7bXjwheH1200xR7dLgUR7cFlHCkkUooI3bUbN1/laCR9ttgIC1/keEF6egZgPSkeKe6+rThwo
ZcvTvS4+K5MOtNqkOzFTM4v5yHLY2xPxnNpjLE153XxxvV80Wg1Kbbux1s6hNf4IgsYcnfRcHMOT
gYTPHnoH1DDPy49bgsO9yDrCB4IJvv0eQ9kS8xQTYYQiSVomm/uh5/LP9S2F0yBCl94xx5icocND
p1SHROBRmaC4upycwtvyCnCg/RZgByvDBXFXcCCzzn9nPpUno1U8JbvREWH4TgOae2ae07wmucfc
pNPkJO1SIGOZm9hwfkaWoDhMTsk57ArmL29BTq6aUXfbhd6Nni21Umoj8vPJYZN7wA+12guqG8QI
3nb8NbgwcwrH7Nb7/ey4xoIbZjP5oUpXWjcbEjpS1PEFmAU/WjXcQFx2lkw5gApdSzfjBppIQphY
jv7FgPJb7WGr4gXqjpXiX4+uO8o2hPBvI1tgG6pY+Jfp55/UcAEnRx8rDDTbAl+1JlJCAPyq4xwN
qTyh1+PSBi/LzigRCwP9h8trMxS/GzQUrDN0LJucMfPADTdx075nH51+c6i9MUJtHa74hnymXRzl
aNdiiDFQ+60Uj02rvczk6TZl27c1KXi7OgraEnSPYiURxH7D0k/uZMfJ2JnvHmbJVrJG30unGdpA
AEv7Wx1LcZmZVmieEXaHt4bM3DUntOjKwEmaN2nUgEId63HBasShjBWwhNk9lAZPnkqhN1JD8CQ9
ea79ZePXG2p68tVrnZKVUR/hoEHRqq+Cr0jZGyJZ3+Fl8guH8v9UN/wg6w9x6lKEB424NTDInvAl
9jv4SkLNxf3ec9Cz9FLn/1B6bFii7j2J8jhZztFTHMiVgyDKhSWSwySLwkd/NFj6GIHDJZUIj0vU
FSJp4kyqkmtUK5NGl22nOYrI/TP3jDSQ1zhTuEXT9NSDdxc1ZZtucXj7tvlgFrR1PzcSAVd0xAO9
xEuiZ3EIwp3lA0LXsW3NjguVwnovB9lsrKwOjuqoZUyW51/U6my/4djhLt2eTpQTpKyFj4ZVuyud
WwpLApD21bMLj9dp9rcbrXEAQ/H7CjpYzjHGC06MrZUtWU3snQ900i3yiTipB2a/q0rjbxmQzvHZ
H4504dHTEzq3WwygZUacFTs32Lp7c2ijrGMk/K0hbJJQEkvkt0Apl1FQ2MlOgkUzUFcya+l+2OuO
vdiv8Fp5JqYFO/YXtw7Dwh8XSkPy5TRrOH37bi3b9rjH7s8oMyUpsyx9BriwF1Dd2p5Mu8RQ98bh
itoXCu2h6pu6+gQXGTpYu7SdgKEEB9kJip2OqYTyjKtJCI0O8a98ntXMPlGhYWTYUJIBeU6a75M0
m0t6y0f0y8+7I3i756I5SNnTD3TbbE8RY7chT9tZrssLedf/0jE7M6EtWYRRc8hizBEIGJRDkqi1
xl7E3FjkkIi2Qji7ClXMNV+qej79/HrmM6kKu6j6iXG7O5iTVG0SyCiFVGq6dwMH96YHWGqe1gb6
mb/ZF/71FNWNzrWJqmUCh4dz7UKkWydtfdg1Jpj9GtrQH4u4HTnNEPnpX5hlKN1KWfYIoHYtp4/i
fyypngGfJOR87epGoToleaqUtx2ov54N0usjNt934fS3u/K9bmdPxPJloSRJ51awu8y9pzsBXkm5
K7FNZRPKIPjCP7ppdLXR7u+xXP+JWjCB/0n+nYcwK42BVgh+nUz3MwMBpyXswuCDxQAQv8DAsgPJ
1cdcXi/6zemcccE4Wi6KRQtjtUFTYbZOSHc4edSpSnQD4g3VgiGI2AaVr7ueGU4F/uFwjDSTNiae
r55NJvmDmXsNXp+DQ2iYGaubiooYW1tqYZYIMjb62nUO0aIteqYTC1KNWdzvkBdMH6XhEzAT4FjB
Fr8aZvBGB5RHs9g0D4HJqBi7q1Lg2QmnIY3XWwqp3rwCVrw2lJsUrBzIJpWX9cElYzITSBPEHe2h
UFbqWU8iSw/sez8S9fOtCDXtzqXgNSxx+Y5nSJjjCWcBPsTLEdLKVzxw5688AIt7qAWrxlnaS2vE
Zr0Ek1DzgqXVpoy517u6l8EKrh35Hfzx4OHkoDT+qnsx/TG6e2gL2TgDTaPTlYR8wwqldsspR9kX
AFqJQst44UomtOJwFu5OYN6TztzyjVK2MzMZz9xBx9Rkgxlg5AmWnxDJ8FlhocueYrCFaNGDiX+g
uf4H5CEnNM9aeKrIL1oz5CsuJBXHojM1w8QJtMiBAVwla09qICElINJShLlau3MJLiDVPd71fXyu
nlyqVDdytA4+ByR/nyLdzrM8BUGLpbC1b77qpUbmfDCCCFn7+j3jtvUanh8/IRaBy89pNpy5HpFO
UxEPwdG6NWhxg+JRT/uTfoZdltAUYxZaJmkd2gnGCI6L5VIfUs2EkuVCG9UnGqHVUbqjUcIIEAXx
3ZAbyGr09roIQljbqDPfxE41xVOQ0RgItHKMgRKRdP9bKKCURe7mYD9qKNodIX4uyf8X7bj3BJY0
AmOdZPENXisCRFtcA7wyMzculv74Bqr05SXkVH4TM6JpSW0na9hOMceCkCdKquuKrCPKQQoLMTPT
+H5vJ9/ktLJ71svMN9Tp4igLHGeL5jv/jrUeItH59W+o5bBb2UvvjaTYpKrNEyxqObkAqYLxZc8R
xnfZhPjRY2x0U7hlMgD/WCOLPUF+jx8JtELYPJ/05SppfuSE1nKw5pEkaddTSRXl0hrnWBUSS+XW
IqIhUSCZiRq19EHImJDUINzcVJ5Tl9mU3bUmi2eqc7ZSC00sKYZ/jzNktGiuZt3iH/CH8OnzNdrX
N7Bb3ksrchAoP0blE3KsEG9tIFFnnbf70t8Ux8JO9RCAkbEbtI1aukDdM/UckPHKy/7JqCx/Isus
wftuIZyjN35WM3K99uXou6AD5QCKaOJGSMP44PbShaZty/7EWlPHBoKJ/0lSqXELT3y9tXZnC7S2
FehUlIGZNc8juFYvh+JPss7JHu5CPbcYGDf1U/CGhc0nNBpSvFZ1KkllqrPVwI/u0wi0n/BLh8qu
Mpwe6ltHeNuhZF28bf1JAY3e5P2R+4GChsf3XCblpeb8U0Q8OOSUDYBnEVqmxUgW7ulZpKu6TbaA
P//+xdEbHk50qKk4NGOMccac0bK31cG2LbqgOMimIpMt/h7s7IJ9x/VGIba0k3bNyUssXe63eDbX
C/jfz0BrLp9fxpXqKGghyfiuIjABYV8WTxEGpKTw1R5oR0FRpRmAulPV9jVkvA1HHw+vVgAoZdec
MZOyGQd0v0kq8toiIwHQamYD8/YreuPXFhvUVyd5uK6J4g8onFETd2Nin61aO5A3kDNzXwnELmCv
OWCfNADyi4zBlrJG+EAMtuKFoXK9maik5Y6Ffq5dwcusWQFv4tDFnyOCiskORBWrORm5+bGkV3iX
AGSVNaiFr1lg/IEENc7pxSOdLBniN3S8T2m4aeqb/AjsALZN1HcpJgf9/uOuMU8qpscJHvWyHDYP
DhsIHFG/JzMOeQWG1P+rHlSnuthdSmmGIzqp0ephYQqSDpoSc+lNn3y11NrfzxVfwaxcglDz1cSE
CAfbWYiFCmWkUgn4W3iyHcMp39rfgx6+WIZ7Zn5/ZoHUk9vi0KUxJIbM8mqRHNDq33qZ7XRnMNVq
dUqpsJKjyW81ZeD1fi0qzVfo/++kTbfzfIiNwGkNAbNGfr/KeKWh2LgWvZLitefKhMhvK0u8399o
iDcqm+ZajLgkowmZrlU7ZaNiSJdE3lT6J9KrNx7FVslsqbXmmfvFx05Gde7cjun+ZAukWOSB0RJz
aKbxJwRCOdVoXq88UUPnI/xMT0TS2L9Ctjh3zRNqJY0sNDLC70JyBURdClTKRsZ1UrzRegAd3ahH
NbUK/3DQMOEM0VJfsU3W3woSkB7cqoC3GMu01y6Pj9VVpwS3Vuft478i44aASZXi3mjm+VUuEkK0
Puj9BzNjsjQbLgtoWFy8KDaqZxxt+TI0O3m/oJWc763uBvG4wk46EDBxv3eK6AF0bkQQLGueFbN1
O0TYviKmYN60pr1Y4AQxQm7U42yKVuPTR3nRlzrDoJQHSICfFToKHySzIP2hQ87sTTnXUqpr0Gji
SmAzD65tLH9CtDJwETnusUprAHf6+bll60SGfuZYNYWXKeX9BXKxxCqAPu/vOo4Ov3uBnNYcep0K
C83L2GwqusTCZfMMAvRNXd6phI/Nn9b50wwBgRWDQzNgF7uudAWtQ6aTn3xvogyhYQP1cF3JSxzA
9rs+ACXNQOLniyAnck/CvaU1Zxye7LDr2sODcyAe58+jzdSHgItQwcRdjXSkgVtV27bYTZgV9BDW
kX5AaA+3E5rnx91vvMzkmovIh1kVOAWncbwYnwclK3v0A85kbrFyYtveLhWgxC1svpX+r1S0PeG/
ICEKuj9O6I8y0PNls1FHh8QrmsgMZZE9KTvxJwHQWsCoPMpvRQEkOWPqtTQ7S/E4GBRjWvcYnOsr
QgUt+JBjPMB9S6FMIOoVoct9T9XvsAPGihzBuB5ZronSvRI6Fri7jNDPk4FeYXTt6fB4j0dwosG7
Wk/naUi8pI9oNJLybD4+sACJJHFlrEjfEEu5YABgvU0WNHx5FJJA9EdafZDMZM/7cjbVyS7RgIgL
kozSvfPxNLESZd0OMroi8jAydu2HVJvUCSj9U7NJ6M9NEdgXinJpKYNsk1N1g1DzTA8SBXT7PAr8
kVfBPrYNo56geqBHcRpUEuRAQiw3X4n4V3wZ+GIfFLZ3dEkSW1x8PknXxwohk6NfNgNUjtcwPXGs
OdDnXIGj3/oIsiU3/DITNq385lZ5y38NQd5AA5RG6mQ2i+Fyy7asTV0SZY+d1mheN3PY6KW9fZJd
SrZH+DHFN2504KCmV1t1QLOS7/x+jql1sGMEh1s6u4MLtwGyL3JhrKzlqPFdUoespBBs/fU/hFGS
Xskba95KX6GKOCLpZ428uBjG7ZQaNX6C+rl8tj7cLSlDE49XaXS0vFwI5KI8xKnof8K1MPbOMc2T
hXK89pCE2+vXnSRxT/Ft3Ivct1PsZO/NMXB75R+2IOZAazVroY6+hTEGUXZnUdUZ4x9ittVRNFcZ
2Yp/3wrPhZnTG+ZSXo2PfhwBrUfk2r8PfJI2q5+8TEf2ofkRfdy+wShnyhyKgMAC44QrvaMdqvri
xXFpmZrjpCoAYAJTNCsDpTlK+nM2IkQIqsPGodoK4goUBCdfLF/1F5kO8hdpfI7oG18ZeVEP9JPc
uZiuZRa6j5UX0RRA5rxqrlF0gly9PmEBYW4rWX6QP1lNAYK7lVxa6YDLWInXo2cuQvd1TplD/WSw
ALlhD4t28CaeysbHqse98imX+FSbbVrWWBjKSWvFQEw7T+EmO9IGhagHIujUQlzHkyS8oFJWPsAd
nhtdOwkGZPo3XluBNq0vprF4EEETrDUG4vEqnsADP/MhmFZQBpAPotEBXiLr8XiZUNsY1kOcePMG
ekbxxp7Ubr9qnuLD1C9brikQrl0oHRTxSI62Mp2U1eX/Qes19e6/4TR4HTbQaKWDK8t6WDqrNaQ4
T8EkNxIbIoMv23BCiU7lzu3xDhF0pZerwrpyth5JI2rSlBQrQHRewJNZaGXh+BwA6+zqxxwJs+m7
hIX4cYOuAZzwtPA7SIfYJny/OOg29JV5o4z3sfCDuPYnunIW5BgUgp6dfAwZW773BWl+VvxtefkP
82s2D+jJeEe55DR2QCUOHtyUtm0ruGegaDJqqmdPOzdRsJZcLBR9AMgXghQFS0FAyv18FWEok9/8
D8gg7AtugmsmqW1fK4eG6X9D9siynFZoT5pwkpRX9CLlknv5XbNhIR1vYj0qgob38I1IR8P4byVu
/GkDvBHi63YLnI3IZuHXz88DEYIZelAxYPIY9h0hQKw7A9be6YLFBXMD3RITMJquE6CRrwOvIISd
j/09DJOBXAPR2NITgMMnyqXIJzeQNzFSp1Y1ug1XckynJ6fTIOZLlXkgOQFBd2ArhukIcdaZUzuA
xcM+3Rb6wKXz+liayLAUgLlNiRhkMfy0AjNQep4XGunZGQuKzG8lPqt/Bgjo1/hIU1s2zX6lHVCh
21esD8H6vrmX3CV9bJShiqDtgbngQ03AmLdA8c5oOdFwkmSv+1uXhXOO33FC+UyA67TboD1wG4/8
qmcyOeX/AQWsMOnNrCmgolPp+D4XbFMFpETiwrKXnbDAxiZJveAruTBqPtX4epE9Qta8t9OXCNBN
0S93BNpncJHxHBxcvkLCRV64KR8Sc6OjWQsly6PQ3YmhY50X/Eod8gBtZPex69rMilOl1UB2HcfZ
+m1hS+/qQPk7yswOx0vuqOn5jkwilpOKd+03uTQ5oGjW13UoKv3phmKmE5NKAMxaeEV2a54TZrP1
0EA5gYCP0IbZVOaKErk6GmkWCnfxECM0eWWzExRQzrI9CQdVshMeAdxXD+Ouo5xkGdyCV4CJmdP6
SlEMXjfe0Blh3RMrddg78y8nyTr+gxwMypb/lZLOueLawj8LOOl8e6JMtjb4GOCyClloA37KFjGT
JL/MhytEJqibkS6mi/AIgDwwOse81mMRUmoASd1MGaTU0FMUA1faC84Bt9MbG3gEUMSHRjqCbx0a
e7OZQKmigZ7Rb7hUedAZ7O7TemQWzkJYQ+jvpK1x6Or6jKpQV8GzEmXDdaN0TlTT0j7QrN0RDzA1
fe0fb7Xo9OxIK/DPZpvSAtwhY9mJOXa83nGfZGzhRaREDXaN2KxR1EH4nBXEcrzECM0xOcTuKPVh
QHH7TAQm7LlcigBGtD44FUmdQrUOiDokc6mICmpoCgLbtrPvkiKLz/BHrlP1KMtXkywL8JMgRP8B
nTrjvEAg/T6edG+zxaKmIfyGvuSIFX5JY1DhruLbM6r6UaxnUzPcQCt+W+BLZ6yoouLZOR+EjXWS
3NEIqVPeYWRso2u2mkVW5fGM2OkMtZlKlkNM0+5fYCyZjAMMURTlu/aQWnue/emomIzYKgZF00zB
+RcxH+toBvJ2PdSriV8WpjupacJ7V8BdvtNo6akPPQ81aZMeWnSrJcKGZsNgfse7cE9rW/Br+vyJ
iLoAGwbtgwz/zv/+nym1gjF5I2Sv5HE4uGlGvbB7ltLI3gf0n/z7jx0dJgXvnmhmJP/w1/GGZelA
2+jPzcoZDNM034XXT52gqhnLGOfghIAhABgkMbtL7+BBCu4F97b9jnRYxVyC14dRkPd7smgwyjxa
mWaJ5q79O6eyIt9+gnEZwBLY7yCiz2MpOInNXCwdgbL2aSwnFZ2DV+JomWKAk6KaAVIG92Jr7uOE
jG8Q4hkZ/6LtvYFKl1Ddzb4yTjCefvFhVIyjaXqsR4sssNdhSXhGIXSCEi/N+oD9Q6AgTKnTtQeW
x9M+8Agk1jR/skmcbCHJsW+GjphHG2AQp9jrTU6Uj/ZI20vLswd1VihKKvN2DlYmr3Qg54bQtibV
I5JssBZ5GyraBsitOM0vw0Rr6ROr+nSAPutvSZB+R7+zD8DNk3TxSzJdCA7NwbbJtP7Drea4XstN
gPGr5FOffWocZHT/UJ7zeull3u0YXWtL7UzI9UgqyFQpynrGNB5hMp5O9pRb5A93TMxdVB3vcV1e
9VJzUbF9WTEg/XTl+yOHfNHEmlOSRM0WucNV5gMzK4M06Vs2ekFU1n+s3IvDRqWMNj2EQLJ3eyaa
E6YyV+o3f8ut12cN590QIUTmj0vMp7ql6GjCYxo3ypk1wmS4PLw4pOSM2gMewAuGMnUFB83g/7JC
nbYZxzY8C2fyaMXhKuw4Pl8LyBpvzp5dANxY0suWg9Bu3OKHIy+Soys3TuQ9b5HxXaghlDTKjbwt
renIaOLW619vEwwlGob3TsXmhjS195lPR1MBbfCsoseq/m0DQufbuvtyYFE0WzuVg5fCL5IPwYBc
QPKBCWoMyUuvjcLuWX4inbXjnhOEALeo+RBZ9GD5newvpnQ6VaA785x6pljamUnVnLrPW/mUOiuZ
pMsUn7B5/qIu6eTU/+Mnsg48oaKGzzYmaVcpxRMVyUnJ+Q2GgyI77dPUjRFjaKOVYlx4BAx4ky1d
2RihrTi/SpBW/ckymbVkH+jTnOjpQLGukvxz1/gkeAW4J/3LKbf/bVlzsrcji2QMAnDu4BARVvSw
Tc5lA6p5mxr2IB9GeY9OmXztVG451T5MXomSSquCmJJCf4t/B2X1TYAxRidZ37rMG+Nbd3kV/RtP
Uy7VDXQAMSPA7chMeDAJl8iLly8Zwac/32R98JV8DYrcPiWRrBGgAV9SyPMO1dgLQoa/xzI42MD8
0RhfH6bhT+3bwCQ1fFdxqBsMnO6UxIR1KL/y+bhCPdg9tQMO8iMLAE4SNH3Qm9yEh7RnvJqttOJM
BWsevc1UcerM7cKGp2uylHQ+7KsFFglDh37onV2gp4tV0K5XRsBlnP8XCLTQKOvVpDL1/24CWkkG
hWNEeXlccAXoBoYqnWyaJ5LsB8/A1jveSs5K/uNTXVi0NhnzDLm/erXywjxSmUR2w40spR4yIj2q
U9IzS6AkJThTDL/09uC9g+MNUEccIYL8mlprbHFdDQHdLpYPNfm0p3QERNpz19Qjrr2NFqyaSfI/
ObYJP8B9huT94p9lqEva60kFW83HCYHqaTgE5VOzzIE06OydwpQCvEhAkIJf7Pb9C6RvPm8oLwow
6iDdWM6AS1jnKChuQ8iMYA1HjYASwrpGdBw/UhlyoAQuef2KgNGv7dQa3AAhkulz9SpEW4Fk0RK4
4Ar0n4s0JeQkXwiY4TgNw2CF1Tp4lXtKw8vRKOc4ENFGjRYgzAtNfHzcc8n/ZlUrtU1etmmsWnTa
xscWvC6BbCrUO8qqHtvcqBVkC0Tuq9dDHiNJPZdIqSksjO0iB/FoTBC7QQmBQ9KK82GqRCViPnWe
/4lC62RBZOFgil+9+wWBinmtI9wQtwCyTdKEUzLjHnERd9K/rFngODzjtoIgG7xxbh8JXwqAPHQf
uaTadrJMwtwPFoJGHRUIS0Y1f3jbg7802Dvos5zBmRtuOGSV49FY0I6vpQrf3yNWS/vbc857ePNF
dZiIM70eZyL27vvvZhHqAPPcgwssb04swmJlnNNN1nBOzEPnq5/iHHlQr6k+ULHQai8JTP3vG7dl
kVSiM4dP964QasGouzO3HIE67CmCr25rIB7wkvVJ+lY8pszA7QTE2g8if9hb6Co7zv1VP0O5wQlm
4cx0faG7lAJSN1tGB5M1IWg3UWB8BhwtTCS1AMOFRuQkAH/Jy8pibVxF4hGgOMHURM7Hg/gfd4/t
Vu4Yc8SXRse3A90mn3pzTEcaY9uGoFF5Yze0mxAxZFEPuOl5683emkA+BHGx6uUGxJmHWpTbp86+
WlDbo04CtRWzDiVL2MyzjLnYaAxa0p3MNI0v1du3kjYKqY2BQLePGydpgktoNYxh58nTnfITgipZ
+qXr2v5wEYvKdvwmq+lwxq0bBaRHdvDtekU/hwX3s9ochLPDgFmmM20qwDWkq6rgO09qRK1NhZhp
8sKBT6p2e3EtMyrZGQWI/9yQMROzBxvUK3UqRPezdPl9X3BZRLau8H1hDz4jJLiSTThKAxhCUueR
1G1FsL2vzCtnTGVNWU6Pygs9J8Ph6/VGFXCzc1SjiT2LHhXDFJGsp7lFdD4RuwyPOXdb2s8uHkGy
24vU2k4/akiAtYR3OOqbXhkGL6YYhso/l1ZDaLpAv4Q1vkHij1WfEkIEFUXMK9Canw7uYs6vvSkW
gDM+WPEegKy3vBH2M026zyGT5JZ6SOrehpCAbbfCgbWlEPGLIkYsnR/SQqLu2wBqA9ovlULTGd3Z
9trSXA1S9AqRTk9xPzKyNDIjGp7g3HjsmQ46d+2RqJUoo0R+mMkYZT4utMLj3hYe0FqaVEaIV5xa
7QiHb82xwzGHay1K4LJR5jbizQ/LuKAph0JA9mPEa14hbDQ8/QFvYp1SAE8YtYO2YaHwv7anp3p2
q8HtchiwncQAqcRdsRkd5r6YG+f+0WuZxxRNAZsP72rgk3OjacOlmLkMgsjqekS7eZjhx+eKNLuW
7x7w0jhwZGNYVwoWA4qAlM54eIk8yn/KmbPHKC+RVPM+8KcMEumc/Wg6XWm9G22q3Xotqn+kGzCX
mkXL1InZsp0zwAFnR5dNVxvYcL++4OkMkgCQfxjlfpedzzNh05swo/p+U2/F87CgNvH4SNYovfiN
oK4C7XkRbT22Xl191+VFMxrGpyIbCos/VZ0gl2qV31lihhpxcYjWcvvFtqpubC9XB7si3o0oMxRw
1Kz665xkHKi5KuKGPtWvtSDwdtY9cwArot8fLITeVziqMsxWLpNrEYUcdEXvTpx0SSJ9ls96M9Ee
sg6AQLeRgfZz2CIGwL7DRtdo9CU7jDRl1bVaphPRTZ2Uz2ir6t+JXTdFrv3A1xycTxqMRKsk5ImD
PIwvJJCUAq84f7FEGOqqiLrdHoc6KKW+kIB8KsSsZp+tPY3CZiifH6JW+2QxCtYqGDoYnS4RE46z
YBzRGsvr9qwNzzaUCF8dzjf5CleYe9/fBNg8BSCdn4ybbw+W8Pvkyn7PV3XHcxzVb8wb3HBQo1dG
B53iRL8Rb//H/4rzaNQY4g5+WoMwa+FrZs66X27ijUpSMLNIzCme1f/w8ORP+lEMDbPWPFvkmajG
KBapm32d7qBctly0aycWgPBPN4veyaZFBtJTMd96GEtUSKavtqoBqw5f468Nk70Tr95RgGzJ4dd9
00TOdNsZODjNNBu+afOeHXNXT+YzvydQv9Ew0HwRuDp6VNUGaFOWtvRBchpi/QJLzg2DcZ06k/3X
blfqDlWPZ/i81i22dLRZn7KTBTJJNNtBrW32ptriqSgOnwXRc1idWOiIfOsMOwfHDmKUgxVzNRty
VjuIRHgV9F5XmZFKtmi8k9LPY+3NSNf0k9vuvBs7CMQpHO0ogjYQ6YFLsO3mWr3QdHReeAyN9FNR
FFkfRODttpPrbl5Rx2X1lmtKbpidIjT9i9y3zQCCJz5Pr6EJFFAKYg+/EpY7KmhgrEDXobx4lO5G
S5+16khwLd9AhZlUJnrFySTwBcNX/e6MMtXgCYWSzn1L+D7qQY+dneB9KyZR35LkJQaur62rPgW0
oaW9rvMJ9rSu/1vs+iZQMnY3AkvWakvIU1ekOjuyNokZx8grOSqlYc7E/RPFf7yIt8VVBXyZcMK7
JXyg5JywLlOCX3PFKs0R7z/mbE27hOeL/oRuqK7jLBsAhE4YYLtw1jX2cHvPKYjnZk3XJ3EC3N1H
1z4lbbNn0ZY9I9q/ZhdfEwlwaxFovkd9H/runExMZlrPAzutaJ/Im3swRPZ8kKcippRKhuN4G4Tr
BZiDJOFLI3dmKfnk1ElwbIx7qcmZaof6FKL2CIFIyq/zC6Vq3tWgNrQYTFN2X068pzAZYz6g2XYC
Ia8UHAxhlsffxn80uiQvY7MvVYuN/f4SwcuJmzNcUn0JiPXY/2GGXtyhkdJm3FEqvc30eqtRJgGg
BLKP8WDGSUlYGn+xKJRriVORTUhB7v6Kl1Dlthp9dWetBLi6Omm1Brf9V+Byj9J7HwdJJVEtR1cf
oMONsOBgQrHBElKup7tb4Ln7S+fXjRJUA8UFXbGZ9OBJ5HzlxAViUg9p0RqNJmu7kwMXm+t4+mDj
yXjaQz1kKtz6Djn6fWwi/2FUm0YLuh3Dmkki6ZzCPlPAilOJ57JAGEPsYJZdc9WcuhbC9F7MLppR
erC0cRQ+yd9r89kEnhGMnWmrDmJBDSCcqj1QeWBjDbLG8D8IZdN3hSzNmubeAAAg2178K+insFbV
LIWDq6G06C9QDN/vA1iE9CwFwkKqkW3jEZRGpZK7XUG1A9sgHLTOJCzjoASalLcRL1pUdnyqF3K8
AsX5gUAC+TF790SjZLhtSQsEkPX8iKD1jFcEYRnv/aYrmEKabpLNB9NwfVEKLPl1vlgzrX94KIX6
y4aUvLaGbAcJ0BuW0Q5EXzobhwBDg58G6cYatk/8+KPCMJ98CPmpejTVSyIy4oqjR6kzLqVJ1N16
3WUCwxUgBmmKBne561n9sty8KSh9a4T45d1ABtvFXI33WhN8/clF+y7Gj4uQ+nKt2EXmIhpKm85W
KMUP+nvfOf33oOgRqf5fpzdeXClNr8e8oMCFzTpIy6mYmIE1DbK5tOEkdnQ8ZiXv87LAglDJlDiD
OR5vXJRqHbrOXItctmzrFkXBbUeBtdJnKnBAR4/cAYfq/iNh7J9SnX+rt3N2j0ZQxS5gPcDxZ08w
cjfDRWIKZ3zf6mBhlDkLFbY8XeP0x9Ji1PAE6zyQxBzXd+uCyrq+3FL6zSQOTRKd9wdwb75uxL+7
ANv27g087ZS6nPIbuMj+zB/QlZiR1nrIUMOFlFBgoG+uzh38jt8VIsBVDvbaKV5rVI6AbzYINXp/
QbaSDzZPuaqva6Njy/Mq4mplAEgNUVweDRb69EZq1k5saY0vdUQUedRX3HwUVGLeoPwVVKtaZTu7
pCwPd8xVxOpofLSaN2bpjsWryUohczxCOM14cryj2UTugsbtFSVYJCx7RFTeYtbWK8UZ/Bm47/XM
QSYOIhGCJrZU1iGmJhh4A+aC+v5gb6PR7Y/0f7M9GHvG+wKXW84TJ5tbTMPK/Vyav9RKmqVPq+um
KP5+t48UCNwUO077ulK7Z4CPQOMnJV6urPizjZagIWJN3wsP+hkzjag8qUOxEviLToF5IZYC6X0L
7qgc1gM/q+8Dz0C0P+zqsUJpA2oG1PftdFXR/zeITSn2DsGd2UzyDKQT21ESEun8vRu3R2SKqARB
XHZRr/y0M/E5jdpqEy3+DHzjd7v6zEpLmPywwRUv2XX7DPbML3K4JMjvC40L2aeYLPP+7EmN7urd
z6b2dCYmpe7RxzqfEal5JqJoArHuRXqPcnDS3ze80Kdbr6Vi2z6lUwuCxARISwWUkbmZ4OhIqcnc
Pk3UyijK0yhQCHj7t54fKhq5J5PozDLKqExreoU+WqammQEQYipZODjcNjp5GJ1VPM+VvHexlXTm
js4gxs4GCT+wgGEJCCQ3XNUodgUkdZICE+rj7zGnUquCEdn7BR1ja9bZmjHmA0XiSglzFHma+HPB
nSx8MTFj2e4cFJXQfsRQcFtDpZ2tutqOCKXBySnyVQzHMzLbxLQ+g4+wx49KhfdR7AroL6p+5XKl
nPiO34VRLHo2sX+BlTk8yoRVi1cgw2sqv6Q3PH64SbRxlNEumLRGQmMTxhziJ+57RDahUa3B3yqw
hDbiKZ9mEpjaFOQKTpeJBcnXhlrtTLR1qPqiJwV6g04SPaTtYhfB96IvO4caw7Bbi+1reVAwomFG
UBKFrvenHVpepDxPK8ahuI8/gB/3+rfsfQI7HYaeBA4XbhUgKLhhIfXkbp9aXllU8RtyC3d2JMqg
WTltJIcizpoC/D0Fr+chCz78nagGEScs0T4EqKmrJnueGLLPD/0XpJzLCJDtCqY+gRsqmQi5usDV
1/++BI6uta1xIzvshTytUET9EL8doyttBWXImjFJO6LQcHvDYYbStzKO6s++iR0JoGC1xkKfkdvw
D1Pb4OCF9PUeonOxhLqid5DeBiZ0n9gJhqmHRbzsVTeDiZQOv+aKsHnGBJ0XrLyRZUBryPRCl6QQ
Nj6YJ8btyt9hBy6cbHtghlk3rSblt7UoSD1n+K/ajjwujKYRSR0ea4VSH4M3exg74vhx6xPK41Bk
d6s1Z/gy+J5um7hG8qPXEjo0XZs9M/nX1i/C2VI5aV5R4NzfMFXaOPKmLA+SBXki3mR5i8N+uL1S
QQEbG1gxdlRUMskVAnx1EE41lQT1XXpnylznfXhStagem63QIUQ6ULyyVpLghCx5hSu19aX2WVY6
hiJ74n9q2y+TNMxIEg9gjn7KaIRnfW3AFiEn78Jc0FFDsKnrl5UM1aOqiKVyhWqwaAhUSZSAmCwk
Ke3ZUv20AD0guZy3hpOFbDrBzvwFFOtN1eZtKZ0VKeJBq9axaWqYHsfDlqMbElCd3EaxaUR5ATSi
DjpgJEsPcCFHAYCV5MlNvsXgAbIGt+7SnmcjQuDFF4mcfxkJ6YHSkHbtPcEDOLPGwgykjtY/iIdI
Qi7s7BDWeoidWG49TNuaUmHRpFqHJbMJCsn104njduXgva/0QSOwCObwS1X3qKV0hJFWnVu+SUsu
mT/cZ2iTmfLLeUeR05h+l3VaxyNYpFp/jk6xbI0i20GSmSrERpilTCzacexQ4mghDFVa30ZMCB4v
NL+s/4zwrMMCRuAQfGSmEm85nRNSEQSNbRtxRLr07jQXgQJNcZ8q7OyP2vNJo1eXj+QnG79Qli3M
eLqVrsSPocF+BANQL1Csx1s1mq5Grxtz+5KDIwPg5AFh18xjT7FGkTMl+aRvVrJFQ2St0h8OrfOo
QrEU3KVOIZx+J8xk3jBN66ERo1Ai6Up7RGQtwtaTHIpcRbhL+pIcXuapjesEEsWTIgtQw4R3+hvu
IVbOUyMrRcfJo78hSTDWhHm4yVXzq7d4hZ0bpJ2hvtEATfetmYogIlMzqI5IpFmRpyyqnvoFtCtf
gS414jJrqE+3B94OJ5WttWbH3s9y+XzNxh0GM57D9CrpvwGfTJ0vkqBMwf7eVG3kuuVCIJSa5q7X
xIGgqCgA9o1VJidLjmMCE+SwEUTy+RDcj1k9EH4h6Go1Bs9d9PkzSyA4zZsH58x0aJ7owEwbWnI9
jfpPXCQpvTSbrweThdc63ZhqxygfeNQ+7TfIN0kPhll2kn30jOErGoXH0YLVpEHhx5CdbWCXAqkb
EPzNGKsW1Lo38Bk4Hoc6kIfLz+z55RrZZHdetYemrHgfsgMK3m7J2Jga3tnOL7oouk/g5TD1Jaiw
qRyDdY7O/JE3aKZHDTZ6lqsX1pbkKzvDhGkDDzGXGXPCyCU4jJqgXGfZcH+xIpMl/JHOpSQ1mFFR
1epLmlMv2IwI4JvS/uj6IpEDanejo+pZL5szj4dKzCfP5gZMsa6Z0g3RqrgUZCCidu2mYJlWfbPu
j7OLX5Y/tRJ6xTD2gtwYDQOuxzpTPH54MRMs0Aj3cTL9ZLkh7DqLScZGTOXbVTk1Go1nuA5+i6Z8
mMr3M90Yu9fXU+v+XBj67PDrPqgamrcmBZFKFwX3aM2gK51rLoITY1wzVwaGiAx+Df7GNkiUfrvn
l+/ZuSXK2hi067MHwsBl+tOHU5L5Sv/KLSs5YtCWNQTvZf5a78JE2Vzmr1PIYDb2pvhdyu9h3NyC
yXv0VVhJ3XdhJih1AdSYncyE5JOGNNtHjWke+8hs93KAUKq5cIQFyFp2vL2tGVJ4/iqftVkBskBk
HjdPlVOQ5DV903r8/Qbwsnl7gVKWFWOzaQ9MWF5u2wskVHN5y5v+xlGga8e/B7Fp+nRw3oSsfHqH
Eky9hTWxhbWAoOYxQliJmx6hVCx39OxeuWbiJkAKUpgGiMJ7imKo3e5+1jfT5PlXCuXmrBuF2mKc
fcomUo7Z8Hl3SDRL+42SLlKaXbfLWT25JX/SF4phZM5WPv6hmDBUJBat72uF5+Ni+vqOKSdVrqkN
4MmFbuQihvaMLOgWms8zSTVY5azB80LzeRBSrb8TXkSKG//uFMdvSXs+VD3BVYXaTA/oJPd1Lv2e
FO3FxZY/oDJfp10Q85W7EDyU4SKjt0g1r7mz2Wcq74s8NWUMDitQjXmks4qy37BkKLKBtB2BTE/N
b4/Jhp1aQQavYW9Oo5Ke35Y2k4VbodZyO/8S1w/Q/hFjpFgUZGDsWWQHhmfAu3onLf6Xt+mQwDWS
eZJjMjVTFuvOKw1VY8yfHVLarwd76GlLxFIbGeKd8AKg6TPlkSvIkvTVYlxsJFiFWeYPR5SD3KNW
wl7Tn0n1PlXkZoGgI4oe61mDNK5QDKsPq/1uIFI4eagliGjxdSmZpSNvD/xjmVWWxYuzQw4B0LD2
smi7SUGmj/Tk13ZX0R172czzmCnZyEuHjKghyZC2ykCtX4uxhGwbZk7gr2FQ6p86nwCcK/odq/Ec
bhIx37+O7R/yTpEt1WhSAk4HR2IrSX7fQXYy75heR2WuYPIGc5b5Y/4W1De2jjy5sYKWqRfyvqMy
1AYnLaeNN3LRzxQOoW2gzEMEVyN7Dveg60Lq7DEVCMoE8NzpuLHH3f8PDAEucKZoeRvh+SsGZyAh
xzXF69vOrL5K/CkglPpvGkl6lW7E/9ETjPreQyKZzpuR6UPXrGeQss1QtfpBK+7nEgaSc0NtdO1y
1+LvE5GAfnHPECESRhQh+2R1SsAZcDBMw0r1S5cBLtD3DBDSJfStllK9ks7R5Cctb/vkqlV4UAe2
8Mi9ZPGPnuFmGwqlcWNjKSnt7N9OL1GIjtYfZwrvggiFvdATOQ5+AWK98KJXPox/7D/a5qjNKDde
BN/OLKADoXgxnIAXWyJ+sk7yqzUgYNthqFoCFO4pWgsMrNO0KGXgferQ1vOfox4OhQ08ixijjGCc
2Lvx1EHAJ2Us0vVfv3qKWh9uQNUK2b71wsD10FICrWwpd8Z871hQ+iEr6X+uUsUsLLofkjSeNQRV
19p57414sfMxKNeT/Rxm4kwGKaF2zSJt0VMmTnU0IHQaeXeu4KRTnTDu3SE2nmQIVt/878ZxIce8
WEpEjpDaVfgRvu3SXf/kz4HWDmdkOxjBtERf+zEfs4lCpwr5OXj42+iaATx/wpwHcn5IuuaqLere
7+iYF+vAnn/HAYilj5HIbaMbXWsnexpV4yqv2KGxJr9qy06RieBr1+PrKW5K4ue3e4Ez12iAC6W2
DkRYNduC3LvvdgeUqFIdyldwV4wkwX3aYh271H5Rlts6LyfHz8GC48bVPr2GbhHREetxc0pddsyU
1C6RJRpAsJFsTIXtHv5EcAQBMH3F5JSZZAOkA3CmG05+H32dra1FQo3Va94l2Wssnb7LJsg0gHPY
gGYME/ZPADQgZ2NOpT04hewcE2OYeHxrgOWOUtPyNKETVgHl03DH2KMBdN4a1zU5HeQgWsA4kx4Z
IYsUgyUBiQRDf8iexZrvjwir4py6GbKHtlwWQJjV8i2jpbk+dlP5mb8rvy+K80SJnEXK6y+iOvv9
4ddtbHYGuLhnzS2AEK4BlOCN2J0Twh7eoifmhYLwSKoGNC+YI7LjpyqO6fb2k2L6ASTb2mtilY9h
VViDlny7dDY/j9CC/2NrF9Nr2UbAK5zKJuwhmISTwZy2nVlAZpNT3NLkxJdd1ukwu4aQgizbGiTS
mzh5OkgkGuOV1zuSekEXB3H09Jpq5DPQygOW35nc+MVb27RUXG3Nd33/k9ey6Km/PMRRxkc7FRWB
MV4g0xbTORZ+AThYGBwNNtUPlLTSBMRHbW6gH/0IBzb39S/1EbcoyjYqQqYJluVJMEKKkI/8CPTl
i512OcFJvupqfJvJSubZMnKwzzg0JVPsN6w0cWZirUXT4mnesQ7QZJeZPE5S2lHt11sbcvYA4FeB
ta5XfBaNVfHCRtqUG7kC5zNHXeov7qPeiUcBc5T10Zwxo9iC1Q0PJ273L3xoQNSi7en69zhc92Ms
SsuUBrH1fzRv0VQ+JjCtd9zOadtC01XXTri/EgBdaW+xOhHIOklTBteLbrhuxsd7pT99mi092ZFE
yqM74HyYP0V8Uh9Oo1Bf++PXF9SkL7m9n2SH2wT+ESUiDWN+Bg3uYuBE7RFVKbEH1YHkTnPtaEYe
tyuiN53fLtCto9+Z3PK3M5cFGAGp74xMbT2HSDtpIVcH/NZYElWMVSxzPNU4FL6uc3fJZz2k6p8C
+eQK7eFjVWO2IQ8yAXg6+IWF5Opzs99abgkr065/tRRXQJyc3x3Zb3D09/HfbtNgzjVr9/6KRtqz
8Wiq9hySTGfqZGoIdIX7ro6CH2dLV9LQwqVvidgzzst2fMyesnIU9PY/6oRPFHCATTOqLy7J9C47
XcAFiCpnURQulQQesIBjd47tLI9FD9NhgvEGtUwK+VN1Zs0T91Mak5vdA93Ytblt74hRcoKliKb4
h0RyYIdXmUo9cYXTFobcBfKf9WyFwketRC/VN/gWm/TjwlxVeyPdOeIskLCYfMmcE3ERXJ3XSvSM
oPZkOaaOZxD9i40KqyeIEqB+PXcCA2PV6CKzN2N0IJTDhLPTExqJqmb4wG5K2iKe3tTnSAcaN5EV
y3fc0XFII9P5DynETjFgCIhRFBLqJbLIaeWbCOoLxBEFqRRzohwxQEFoswXP3fMlQ0Ovvta2yQKQ
IlqjmHtWw7l//v/f0cM4oNcwRJUk9AdecpqiAkT5jEE7o5shcA8wiMAZrUAwm1Lk7bqxc+IR8S5i
OAFYXpmtviZExc2HdfvQwV1Vd7jqULw8C8FEr/G/988SPgtMmv5kvy0Svf5DxfWPH9mPhnKllDMr
ew7/zPZOuTzc2QeLYFXDAmPQn0ap3EQCRNOw2JPBEwLrdOmGiLtqpJCVhTb2lc29rGn1IHUBxtsy
riyaCk/P/Uk2Dbrh50NVPihUV8AZM35yCwiOe+ryNgADQ2zkZ8mBqPqqzWGo3WXg1xd5O0fAChNA
tzH6Rn7CiYlxmx/vHQqQJz9X87NCTsvr4Xxppdlnp9E19DkWBN/p3Cc02RmG8yvO6nWHhU/QXu8O
OmCcxgYfG/BiYT0kjGIdO0DSQwZQvbldZ/HBQnOnSGhx3+ueQPZx5gn6DNGRNijk8zgYnq1w3VXs
yQ0ORoxbhhk50wLBzSL67FGIkOYxn/GD9ar1EvUbldZ8LgPhXhx4yBaUeH6qr+mO+/mhR1LfBGyW
A70LCCG1QLKRmBK4HyRyEYPSTW6HMvSEzr7BmMLqgl9L1svEnf76ZdluOZiu0Rvsykwco5Kh5n1O
2aY7dtXUpDQdhqNgUsTPfQy+SzXBjUnGJgLKvNLsVFTMGb54mpye5tOqduBSSWdSGSF1pY1KR3+K
377j5LtHT8ta35yLRTzOYetijwxg/hxhiBH5dfvE3GEEhdHj7O7hHpdMId99uQUzSZZniQB2Kso4
PzbBroW4cu0lrqSHEdhpyspGi+B477XOtKopfpYdCi105ZyERvPGEqowQtuckG06mRbaU+KZBi1U
CtYWdNfl3Wt4ZFARLl94Rbq2t0macM/dTGJnT4gEzyZGqvd/d48dyvqkEBliEYih7AyoV2pnepA8
vf15ogyBUQA0/lAYuXPz+5JHHCezikiTzNDoEp+HZZA0ygMbuUtcq/rsuGMMkzsTv7y2vm2yuZZf
zEHA7XgRDppQALVVZh+qrbR/ovz9IMrCcrsOT6oz9fuyjpWxqxTiwpGuIqEv8fxZxgcxEOYKaaBv
bIfuYQOoJwEbpG5tuQy6LfRm6SIOf5Rq0/3TfQTdwfIm3IxunbX+cmSyAOFQ7vbdw3HclNNEruO+
EHmCUF87R0WpxMN7PpSY7hnAh2DqwsDT0VcZbtT6mHx7fOO++RdortAgNOodseJmUIgbrY0gdoQX
6UFC2LnHnWWXqZ5Mv4npu0Z/yT1IBnuxFz6eAqoMbMm3tvIMVyNKrV+VxqdAO+7RN4OazQHvD8gN
+rb+ANzx4JtLWbsVeFq0Fa8IokV7QyNwEqeb/xlZNa78DS4U7niZXt/uZ4FXEFRc/jil/0JsP2ki
EGI1yFBmYnETNx5/J7UpAYCF1WWIoF7BPi/keF0d6TbFbHCOnnJ2zPHK17LPNuPRa3nTP/BcAegG
HyiGgdOhLISbIMnyeyBw9eljKklPFLGm7FwFa79EbVS/DYH5Ay1JDK9xu1x6NXluCpFTGfhq4iWm
jhscC/UQvoZkw1n4F713bfGztJ3r73L5b6F37+ZWoE5iPmo0UrpXVwqFR2vikPedTNvYfBRedNb4
EeD6blrpqj0iSx3sAkA1VoKWqm4jBK129MCWYt92JGr7tOkw69rc+thun5NUgAJJLBRLKqUIAFth
NjeCVDw0fsEsV84EW4bZdojZ8Yzeb9DXmEqPozNBj2o7WZggi3osVmE2GL8PaguyfYThYKbpVa/l
HtZAK6E2X53tkbtIKjkdxj1xnOP39JVpZS/Kj86RJC2cpgGwwRQ4vN8K3bALWysdzZWkPocaC8aW
jMf45g/GwDggR0a5KCnvuPkFJWG6EjMH1/P9/Q2yXOH/Ar2UL8Gc11gEal4X/teXHyTz4NXsnLSy
kvxZHON4MJMZISmBdZRv/uZeAf6RvQFm0XnmtPsg6G+Io8PMnsM1q9nYqv9ndpQ8vKYxPEhRq7ha
0o+a2oRT6YLwCxYcjjat1LUCiMn28Dvd57fhRwL1jbPWOEcPKiPp8JYKMQN3AAg+40hByyAwLYPi
0nQQ19iu2vij2zBXSiWyymHnrfsEkrGzzw6EWJppDAewFlC6eds7xIQMXHSVOnHsV6gOJXjncpe0
tTAi6LKLxqamQamn36EIFrFokHZVxHnsY4Mjn9A8+fPAqTZ8XzxA4byCPirunGxWFv5BRmMY6SCe
fjXx2Y50FhwF7ykf+qp+Owo5P4w5+TjUTzggf4FYPFwbkM3A/jV0G9evGavsd9dew3rnstkGuXbM
Ij7aXjULwjRPA/DAzfH2Jvmh8cN1DyU2Ymf3FmZoCHD2hro+SzyNelP+rBKBVhluQflSlfFQwmjY
KCAroVyQJaUcRAxT98su1NwrwUkPAMCnEoezHCW2Yjo+vMWbXLGZ+33zZ9Hh54xXeN0HSmsEwsGs
v8iU5mK4zNBhfuUY4RhNK7UcsF4N9kAXJVwBiTGQ4XIXkQeZAjJlLy1XyS8fSi1f7r46VqyB49Gz
tsw3Brl6q7v8mu2Dy8J2JdY2d0I7zZp4XFsVSUONBoKmF/D7bADJlB3ykr/Nr6zkGUP14ontozoQ
AVdJF2CAwAEcQ3trV+XEls3AOdoTXd+00GdAO4ybgOI7Dga7i5jbqhqMDX94+2CI21Wb+IA7wR4D
8WkgxM4h+W2c7+a8kDKMNiNAWOtnDW8DPPJqOB/1f9o1idQROnRHc1FYKNpdQId2LNPHQ4kyqO0D
5zV2SfpVnGWW35EbV9Ea7nhKpVXwTN3XtFOP7bi8D4QE/SO/9B+e+dtDqPNErcFJZPApNroqbBv4
WiTqmui6XliSLzStPjk/yYafLhs3lnKZ5Xu12bplGyNJHuUbmM2NMx6fMDv+Lpl5ECKs3r7Lb1K+
2/e9dSIuhg7jqw2dRJYv4R86Aala3WDDirTGeXd9OhYfBuSiGewOPh4sSzLkYu3dpFE2XvfHSMFd
uiMLPRpny+1TtCjFja9kX5WOHBWab/hawnWaEBErjRr6i7t8Skzhs9iBKMGIgxynjpAY8YFduwWM
fYr5jlBRhPsyHuiPl3FqDO0NBdZh6Gvo9hYVGbTaiSRKNL/oyorTFZJvW2doz+L9DKpYXO4WfVY5
G9zCfVZuSj2vX70owy1ceVSrJryQiTG4zmcu4SkfJnkLVuuDv5fxQPse8KGiuC7as8nnvdx/YX4n
oaqsI4EMtXQL1GSnp8W4vYjx/4M8D0A9Vlk2Akkksxx21gWSB8ltGuvQaF3SFPYCKOW/xyQC38I1
9nryYym0UgeVv07DdvdglEo5weC6XN2e0yW2Z6MQmIIZZN0Ua8HlsKeN6hHEfNWbI6Hx59M4ENrZ
RxiiQZQBUm1DO5SuoQCk6jRDMS6W305+oQrN8MCDDbAUi6U8NyNlAXXR3Dx5lpdE7vTKDv6MFAbB
yFttST5IgZ5E4qijEtochrwwPFbvgnyfj/v2xIe04d8eAA/dfFMLEbHuabBeFv2F/D/Hp3dlmNil
qiojzxheTfcJ+SDfjjVlcpjfaDkgA1lP48dsRba5XraJhG1Ki/hgAtq4U17fcrNqkKvxqEHLpsoG
hmA3NrcB8QjrtVA0Dqv9jl5imClXCQPwA4B4Il+azGQ5YOPrDXg5iyiMZVfASIiizzN8yA8uWRbb
muprIDfwfFaocWpQYUt5F7W5YaudeTy9/lJBkUjp7U1+uTVyh7Nbwapwju5MMZ2Ievu9+Xrlkpvj
GxePOwdwhlFwTGaz6cGr4oXSxwPbVOsaZtzDOijqtaZPT6iX6LdlLE8DaUnU8wpicMoGc8Y+Sfbx
TMKCK+PEdRIRESCCUq0pmQp6U1l5/o4UjILsYqlKbABa/+kRd8D9tlzsrGix16mJaRvlipRofMlL
vXDCU3Yw0n3KDOSnpTPKOvqb1HzBSHXuZnTa+ZCKo4o3EhEFtjy0xdbZgnM1zxWI86BIlf3GqnEH
MwNbu5bkpABgS82ubVHqRGF8xmXBNOrgJq5MQeLEh4v5o/V9gspcgxbIPXtHccVfcapMWlh1hGjk
DUl3VEdZXxjIYmYe3KtLCIjzsWDw1u37Y+wya4gInzz32ogkAxFy3du5kcv0Q+lvQWAmU9zjkPeT
YLdW9hNj25FHyWHkElzpTVc44IWVqVSnGRo3FCWDtNETt1t6dM94lZDZnKuf0yVh0OkzJEIJ+HOG
O3tMSTOsnfIoPqVAqA3D1F7JLIm9h9GHRk22aPJHKAUdOgF/oQdrxySMkKRVFR+kN3fv9OqAfK/N
tndR5WlFgT8e0H8lxYTAhXd0W/2Zr5O+MlnquEx4cKVPOKDUOfBkpMUdhNiKqMW+7E8CwB/UnnjW
PVKSsOjPal5wgSC7GXkKZml0EqdhdXeG8OeJGLCqRfb5MEyILNNm1KO6SivytM2tu9UkD3nc0sQP
DVaj/KEw+3oOq9VjtP0y1hSxIZaX0QKL/6w8/Pb72m/helqng0QaXJFm7VqL8y5N5OmS5KwuYJvj
gEZZpLbM20/JUt/mIyJQzNf37rpH3j1sOUKvs/PyZcLownsMuTBW1p8JC9XnTX4gEEp/qquVjVz+
BGr3t6zm1NfBVcuIgFk+T9yv3vZcBluRg5ZEzRehnwLccNvgKxYGM2o8azOmdU6mL6yowQBZbWQP
xVck4uRR5LkI4E7yNynLpQwVrluV+Nfi/BEdYv7RHIYY5o9kjAxSV/y50nn5q2Gn5vtoVIbSLuEp
Edj1HwHF5/3V0n3A5GE0DPsePyCpTXOKk9nm74BdAzDH+a7gkIf1AsMpNPY05huoE5IKKZV1ePzT
+3k2Pk8+G3nBWGdhY5i0PR4FW1BPquqj/Z/sH22ImBcn2+u3xnTS20wCIyuzor3jX/EOBUTFqrir
Q5FFc+0NqSqNxmVNuhFdT6ix30VYHDzHwdSfRZBi788VWwpmQu9VyKcbzcyU1EYUwAWS1bbmhKfE
HYsy7VaPzSxRyENjZlfaP3yRJ2//1RV1WfXj81ud80NdjO26sC+qraY8EczsYEcYLBFY16cLtSHz
uqBAy0tSs+q6tSB8lB4vKEX4tC0a6B/zWRklIjOkbsey1ygmY32plkJ6YUjUeF0fHmM+jBm+z4Ge
Hn3XQ2Cpoomuwyh7DK4ODTFceQAbGDpSH+WBfN6w4ACAaKJiVFLcc87huo2MKT180ZiZNyIyFuk4
FePbNvpB9scbipIFckIg0aGmxsYzr+39L5oppSj/bSkkVWI9TijiPHlR2RgCJG6je7jNoj7HLg9L
vVTuEImIiCWYh4RVIlxLxzNQ1apiUqYzg9e7AJ/rvs4FyVCEZS9jVyNB925IfhLRAusH+BPKOojx
GduFBjYTvq4W0XHWCDvxY83MIV7W4UyUvIvqzTGyLTZNpusaCKsU1pfFRRUuSAZTycmnO4JaQADB
c6Bn/B9SDz6Vs/Ghr0QcSYNkFY1qFHN0YrEHdxJcS3BrDh+/k3wVnVP4EalEyXc/lbD/1hRgCp2P
jsLzbf7YxpCC+BdazhE60P4M6jZcw3XTxBHbTO0cvWogZxh/kfDWxXfRNxR5r7CDBT6IjChUftJb
NJGMhxa4kxnh+ZvkivSRmTj2rqDuotkw3nhtLLKWmtKjUgEk15YKp9wZ/cVZNQ/HWVUPMIyYgZTe
pkqS6Ioe26979ZwYieIEwXH8gccfQAlEIpSVSjyms25vFSwutxKp4RRg4mp8ABK/cKKsYtjKQhod
M+F91zAiGtsXQnFTfG/zTqdZOu7fovj6U8h7kFgihCmY48EZbkysBhMSAgQzGwwP5JA8I3ZL3xx4
LwScG76rNJNgSbhPP80N3dUD9OZfqfFB3dwoSzczFRJZgAPA/FNbfXQD1VkL7t/nmXTLe8ZD/4kp
RIOn4hJNuWIWcIFltq4TawXbTw8bKSVsHDtsVaAJqmeePILi4pneBwRZD+/8bDo4Jlp6UYC6KXdh
WQDQIx7XXrcTsrB2Cu1c8izfXkeDK1xmwsTDZrxi1IGolXs1B7xxpEHvjAGg3TLbsfNXHuVnPZOA
EPdkTaKIDHfwnO9qx3QDiV1AHuGvguHq6Fc9plv5pT0zRuFEzRe1v5/KwppFRjNEsSOljWuKtCEd
exGc0+9CZMNOdXOHxgPzRVDpTQNOdpPUgLYwaJdLvn0o7GAH2ycRQK45+a0XCs6sHaXRo8dPqbLX
ZrJkK4xy9n4kA4NwIqm98lVVRKxfJRLH1777014O0Jmd4D/qMYCqU7LitOpj8F8NByGEt4YvJV6E
CogluhljI8HvhdM9lGlpcPfh4DnK7YTLuvUzqiRKRIVHJA/CujCTH1eLfr2WEXharP2i8fkKdtlK
O1sNzvZy0tO9VDKJv0dBn0yd0tR2Gek8o57bwGNFEJuFqPLre7FRW/4lXBnCcRqwLZC5NaWUNLis
sm6O2hpAQJm8ksJum1u6c7uRnd/wMk3l8TA96eazhqmcJ7LGyE2my/0krJ3azaa+zv391/VmP9vN
+C2Tq3JHWjh/Dc1aABcFgUDiANMYXgpn324NI3LXalJEIYV09NsSZu7+K2R0JLDauY9u65Sk1djg
+45lcljQi9hFp90Qc93ha9W6qmvhvig6MkPMSgJZFYpFIMOVhCOXptkQc2VTWEOj6PzQQCodR2T5
wWyIRgFpWh4p2xMVFcVJZDQvFbMkCBkrz6vsoMNXQ73N2Z87Gq1CskoQDKpuggBf2/7XgxzB8Qjk
cGDNbiQpq7a10uBH7jjP6pPrKtaO0/+zjafWePwx/0WU1rzzdo512N8BFuTe1AL3b9q24bibzjkf
e5BzzjspejIq+sq+5WpJj6PK94vaAyyLsB9HyGqgF+fjS0ISXRlheyR1a5sjk3MEfSmoPSY0AW3O
GMptmYxbMK8yVF0S4N7e5ROXhewy8ET1vL1wi0hBQF7kHagSCT2X18qNBzZbFEhxj6u1gwqJyAAz
vSIJyNY97GHQJWL0V+unY3sVh2DoVLltN0W66tl9kb2pz7TsOyePG54D2N3VCT2nHbcS5TGekOtQ
RLLOFGAMGZ77Y19ZCco8tExJ42F/zckAQocEr724yJXzoQPhKN/n9jgkqVJeFXUbtTe4I9L/DpJi
bcHuRm+W7O4RfB1K/sgsgsup+Q1dZijNukit2VduB3nXfkdaUVA+D0OPyWbSxY8wq3ZN9XQyymeV
TV2d345OmyAr9rpa5FLfZ72rQqhygWavmSHeO0WU+ioLJxxvkE6MY6yhSWzIEzSnULH6RFvRbqL8
p2KGt+nvB0RBGuaTpT9gQ1WSy4LGFCBNZ7eSwHfXhUNBJekUH+TfnCHF55hvK5BOYugrghrul4Md
iUqLKiVPX/JusT2imIu/b4TgPHJdhdJPj23SZ6I/8TrV9Tkby5zLZPbIGlIDMbkcCqWBDRuwgzaZ
uuIqlUmmctkbZpsbuHSqHAsZlZ1MXEV5UTG3oYsKw8Yt2s+tkNtgUb1MYZRVVyI5AEzZ0/KKCpVt
VJv+uEYGSD4OrUpCpJ6V5VSbFyAoC8Z60qij41tM6MDT0X8RRNRKHLnoO5oOYRKLpURFvc8tCwm/
aC3hJ/disbfZsTf4W3NPRHBVzozh5aLS+r4KdU4Ot3VN7JVaIUl4D4qm0S5LVzhYMRJg3llo92Qw
PVHCIiUnX58dBo5z/7cAVlpJfPc5ZIkh2TKiMkibfMzqo8OyAmwZewNa3p9nQygg3jpjyRl72M+K
c+d2ASSdz3nd33JK9LsQHno2q+ru9oOA29stp5+2XqLHKUhDgL4yNREiBiApd+wiCcWOsg+kLCBK
KdHiwcf3L+LNiXjWzRx1Jd01pR3X2XmKd5u/Jc5xtXAk9TYfnKOGksw+Tuc8VYOOi3kATu8Db2ym
53+Kl1D3cPTp4bqlSC+t2YlP10eFbTxH2uNN2XMqzhYOnV3CyQ7IjbptyNlkP1zRDv5Ai+Fx5qDM
6vahWvkZrjxDGXW5A4zbDIGHfvJsrhvzajxUeA3tIPs/9cyQeIRQG/GZrm3qCQkSRSSii2GZ1OFO
Jw/r4IaQN2FBRLe3qCwZT1QYlly8SyjvV3mf1WYe8jraqOqxePKgCwxf6AXaccyZdkRCc9pMf2nd
/LifK4bY94ZiEPujXoEOtV28s/4RVASEFJ1qjy2haX7hTqjUqzyPMcNMBx9+N8KUi5pIh8cl68UT
lNwCmjUdSg2BAmIHfGSMHURTwamDDqWFJwtSf+E7yb2V4LgievRX43kODxPh1wmaYTW9r6KroYEk
ENkWMx9XKk3gzcwmgqDr6fFzLMuKXfHFJJA/S5et8dh7HKS/58LcaVXD0PM9LJ4KPR+e8zo2mctE
FNT5KvOptU29RzyK+yZb8YP4SiKIyPrDclcYhrMoPnE93BrV0ji81wGJIu/B+4bmNNbx1tYHooPo
riO7l5fHFihTW54kSL/tc4XeOKYvovyumm0SA6w+MH6w2SdRWzbdcH/Xgm8HIAd5Bt2lK5/6Tj9w
YFs/KuyebopJKCHmKOHtWwInEdwltj9pMIj8zt4y6Hgwcm5vD/IO4U40gefmythTAu0463N4xd0W
l3ORT2gm1+JTEn2oLsFOmwoEkyPOc5zo9gvNMXxM9BDOgxGrJRnzCoSZU3SYmIOlP6D90yanI5/Y
ByCmSm0/Ozup6SG64mSn61gOk+hSRLKqyb7F33eja+xBmdTeSxLumDK83YunUi2MzxrvvZBsOqdl
6LfNQR4l3db/SgE5vn1rjKy4bhlTHYwOfejdPhr8mURQG1BnE7LS1GNdY3297OqccyBfRqcgRh5i
co620PbLv5GO7p/02gSmeL7N3wvBqxFo7BfWkKzU1QrpL8qv+Jh/93l1H1ZS0JYFXuvbyZYh8oB9
ES2eujAVImSoftsSecHvpdagkdnxIFAUyQ28+hZ5Z96vxHIW42yG3XjKVbHZWKqGLdPNRn4qYl9e
5ECXBuUIxEFQ5UwRrOYlFgUjq3c7M7n0fyFNypuQTxMrwo37A5R62X+/5J1eaJQA8XV8rAQbqLMl
ENtBOzoualCGpe+GrYjkQPffUuaObf8HcUWUkTf96Yfmt9CJGRRS/A2/rcIQF0uEglfyNdg/glc3
R4evL2Ogx++nzcajbyNL56fQTB9U8ywOFNOGuBWass6iQlPVFXAr2OPViguMtbWWngEg/6CEk/yx
t+PwFoTJTcSbOKg+NUDjtXrUYqDwzeVuH5CovniKPU5yp7+xIT7oLL+EZIbI7BK7LyltrZ74K4HY
jeT5pqFoZzQK+w1nclrsvnhVPlgdQ7MY7LcV7iaGY5uT9ph59NDIP59T2spEXv82wKhStA3JOesU
9QsyvXKTi2mONN1+SEPnWveTFRzWaEpnT61/xYwdcCK08Vi9EdX3K6CYKqzK9gQFwZEbGzzcbc6C
FCfTRwfKGZlYFjl5K7KOM01tW2xz5EnGri9FgtC0Smy5BwydrXA8mFIXZbtGkXeYbP9G+1hAdPDY
83u088j3YFq7ydjLhcwd0qjk74SyR5LqFMJ+uTLYLZmlcuJg0Ry1iTJGKeuMMZLJAvmGD852ztYE
VDjy8bA7m2gkw4XoDoxxQDrFrICL3sttxo9qf63tDq9cm4GAKUncZNd1igA6cjniEbfaSBWWxPZe
eXFFY1MJeu+Cr+shkkH2iQgDPMg8kAGFeBg1TrVvwcIpP075lGnwlLIegZgNmZpz6KYWFO6X4qa9
SfbxZrajkJGqPgPLSr0GB130jiP4PZy03VLbGkD30GFcBeyHEmG6ZwCGR3Ltt8Rq0ZH00XGZm6cF
gtHtFtLSxhCR8l6dBdZDC/qxo4yLJp4w25SU9OI2f8Lul08d+XwAfdPQf7L4IFVjeCUDGsheI7gw
zN108sXKfxc1KPnP+8I1cemf/6CMNxUiA+I8B0sN5xs0W/or7UuoZknOWYORArvXlENuJgcSEZh2
9QtVKT0nnEVq4h7bXxCO8F2IuBCE12GDVpGbS03KwQ+khm0pzhBXw/DM3C6Au8pMVJ6H4fmGTAC8
KBjSA+VOOvKR01MyJBCEJZkI65sbeqDcM5BfviN2XxXNbRRlD4qlsjp6j82EBhYLBcRVdCHhKlr8
3djt/DJCwmIk7Em5jgXrgaXnywWoUU+iPX7SGq5IqN70wQZCuy0RJEzlQOOYmqk1YPLvu3V2kJLX
jUgfIWZLsL1Th+0GNskUfG0CmJH8/tyvd45PlGOTk+zgaCJSuEgAQUCtA25qIXymyVe9JlSho6kc
LCXQOjkTJzVDdwRSX7Tyw2QpVu+NGxhovgGIw5f7pfBuA3SJd+lXwyd22j0GRLKJM+YToDwn6w7n
dr3bMcAGVz3UXILA0+GF0vV+SiaUtMtOj3PbGTKnlG6HgF2wv0ljQcO0dHQaeseWoGj6N1eswydm
IqCoZKFVjsmKlVSCWVlQl5N9KNslKweCQ/3lLauzL6hkKL9t1j3zBHq3kuVSgvLKcs2CHlRjUgrc
DssQKAWPpBLug/A/Yt8EU5wTQo6uSz413KDCJg3zeArI3PKL1K88Jmb4c1keUxaBd4OrsouOePbX
rxqztT79Ghj/d1l4oZYkGw8Aw8Z528DmK+B/rHOSYxzEL9kU/LpYeq3Ivtad4q9Jq6gfsxldPUn0
EUoZayJrkYvJZc4cXu/7V4l4+6Ef5/MeFXp1s+ZY+7ucdAtfQS9lHuEk8C7g4pyVRJ1xZ47ae2UG
8e7nRRZ91ZRLT0GomYwII4XimD9PqnLUq3YqEEmCtl7f0yG0Xu4hQC8lSdktRJiHpdQiD2Gqf51q
YZLwDYJBlFQZyBnbTXSMiD+UtdGcHgQr/PXKqA2TG3RY6PgTSy9F2MZQJSD4EdnQ9bauNstQuYa2
6iv3AHolJThNGmqdO/TamhabguZkmxIz3QC0Za87Tx8LHoDOTaNNKViRv7z/glphUK9Fg2hjaMyo
ziqgmEbbXjpGVqLDsdFURFxblPpt1eG4ZFqtyQ7Dd8ZQjqfLErWhSimCUxMB3YdF+yBInq6xbjlM
NfhLmWteUT/8ag57eLtCkadp40QDW041+9Q5Ha2jozcge8WnTacghGgF3mf76OJ571cRIwCxfp0p
K0mulTwjWQICi6i/623qnu7hfwjuJNLuoouYc+CQkdLzBQcxTIihhaKYyZGcpHp+wQ+3oFKnFGno
9P3VNUv/JpHVAg6i6gGpjPWBibg8OuWsvk5Lv74+ixnuHTQ9WK8s0s/r94GbS83LIjNBSpHWOAzw
MU9Z8VkDS/Jx0ARl6YJs7V9WblNeEbNXk8aqfKfKJFfXmhNCg0ZPWdII48yZyqpflmmNOI6Nc6KV
J/ZpULr1GNdf3dK4RzUaWYvf0XT8K/zVUFi6xNdM3EU/MwkcYBdwjliscyZFi+4DGNYW6EcAMlFT
gJMgbsjdEagWUokwVgJz/Lyfudq1PyhfVGTCEUCNxq5q+OMgnSW+Kn7adkO0CFzWSt+Kgs8OqSHn
WprZq7C6S7YCWlh+JLtLal4OdLwsd3+jCj1s6v83BdYavXBHixcmCbWu67grXOZfeezp8A0hZWcl
6mDj+62F2PLrfvNzMddfLb9QiIKQwELIYq+LIC7rbREWvqmhDpzYy2jd6ZdmiYWeQ35RkQP4G6DL
pZdxggjE/zzwNmOAPnbwdzRvmJJ9V2VDi5UChIDuGGAx2Fcva68LUCO4srpCYhBjOWXvmsN2FKzx
stD68ci+HROs9LGj1q4a1d1Tib2WStpZs409zPvaTxA+7YfnI2/s3m3ERVMDpqj4w2FMFgyt/M6l
sNG7s6OG4YWf9rUkxZGUgGkbqm7RDn+vhsNMA+OKC4mtrTBk7+0ZBRWJjL5JcV0xQmUhU2lx+87Y
coPNp3N3fM+tm4nyOU1fXc7O2soXPdXDXnFJRCVaHdWQ3vtWX2LBcpALU/9sliEyKJwf2KUcsybB
wf0xvwoI/mbk3ZKqL3zeHKC9izHUZZFSy/yUS8OVB4dw/OlPBDOSPJfeyUELyWuiDEKsY84vz9kN
coYxAcOUfBPyaHomdW8GpGih5RUq18h5eiuNJUjKByUdT0A8Zb2NtOH8dMZlLR4WAw7sFST9zlDo
KJDA0w0XFEivTZ+mZvkiTd1SjjHLIMRGdkVSZ3wwZowSHTskdhNs5OzdwpUoOYB1ytobQkJPmixR
qRoAlwpeiBEW8RH1kTpto+c0gs3bl3xUDQuh3EbSAg4GpzJibz9JdvoHkMu92BNl46tlotjznlwp
21CdoKsXxr88LqVhnDJ45ezqUyEoSPrX/5DFsBna+JTTo4iwzqi4XaYGiRK+tCl8JqVxb8mNLMdH
KKcne4hEXNViFb4toU+o7RAV/Cbl0fjRc1YX8frVVrpOP2FhLBIBRFpOirVKyXlb5vLQi8o+dPC1
2oUus6XHrsCZ/iGQQ3DPN91dZ07fQJTe678GOk24J7fkvlRhT9ppUiwSxBOnZug6vTeFy+JQ5Mlm
W8K0P+h/NqlbTaphHQHes+iaANWgqiHsJMU3YFh2B44Ey4XPd4YGq0ZtS+pnn/NtU6XSck/ZXWqf
hBYC1kyTos+pkP3rYf3Gyn7v7mRXqhpkgwnDYKfYleHf9hibBPOGDuJ4PLzbAiTD8nb7z90NmXeZ
LYO9f3rUSXvsYdogL6qh2wXS3Hq8MYWWXpSZvalnU/vfsejbXsHG1cUYxT93+rsltfVISTiEX9ec
dy+KZNihA4OU+nH3AwqfqLGpEeYkX4s3rT+JginGtW6/WhAzSdTEaAF6ts5gqtnQmEX405x0iDZ7
4Z2GVFqqlUAWLJCSEbcD+7VABnM0ax39i2xwGFr0K0Rc3OSdDm6KstW6s/SUv1TxoICPi6LyqnH/
s6bo1tij1RkiqLwsN6W58N19Uzr1vvzCiL8/RsvCtkBg6MdGwXnOqEiBJ9fvornbjw5Zfpe+3mX2
sSh1Zsc8o+98/oyX/2JWSOBjNk85leLG5QYpl6gUIpP9uGVGGJa/wcOlS0ht4XJLtqLOPNgI0iBN
aMzPfA496JfDfnY93SQEHiQT4PfJ9EkN5yyKc75/yuqBwCPmBp5CkcZ2ihbCPqwjd/mHvIgoN2m5
MPJtibS5mJfY6PypgOSftO+F6bEtN4nLh79Hvxv01ZLvigfnhjQ4EsDnFIfV3Bgaymqepqi15s29
v4u8feGle10bxFRYefuu0nc4ivVPJK3QIK83BHfZJ/VvwwD3al0ydF6/qwbfaLyHSpfk0Zvc5SNT
L2QFnmTopjLLNTmd5P/r39RGbu38HVvpGF7qNbLGbcPFSWO2JAtkeZ69pRfAyKfC33xceYiJDxBR
fMIFC60PJvbWhXRMeElZ9SjMg1qHmKLaOaP/muwIH6ySk53HbxE55X3f2WObgzHxv8m1T8I44jcH
Ib5QCj4Fx0Q6/QTbfDHCgZ4DzwXH/Uggqm1glNg1xG4kEunKqAH5VOUKbmjTmW/mfOkYKOPPnxnf
HYrx9j2ncnEcHdbWCB1sJX4RQ6G+Z/g1WZ3IcqmTBapG5m7bD1o1KsexQXaleP886D1nwgsW/VuZ
Dgcf7bbzelgiEs6BDJ55qyCbQfrM6HFJmoLConFP1kur98UVGbOuKvEgwBQXYZibI4hcJkigVTOf
fuGl4in4LcPUm4G1hoS1SH7Z08S6G1nri4JO7vhrYdd0HFEsTF/i/KUhht1Yij4k2orTy18gap29
PrBggey91vz9GeqPifLg1LEbNajJFUl0aq+LlzoA+oNwz0VYQcXGsLasCwPcp8OGpZ0ETfgUUPqM
tXBtWq6wdQuoIlL4b7ZJCINs1oFTDQ5imBgatX3pn5tOfGhrD+Ln1+sCA0EL46oR7A8c8v4USLkW
icyTwB0zVhx+D+D1HFqRDjK1jAS8NVCDNHfgAOaH4diWCA15B6Kv9dSR88EkaYO4tXNGHbiL18Lk
GFtTPYQEqNEMNWn+/pajD4g27HNlXwFiCgubjz3D/07ejOWzNgqqB9wS1mh93FjZg2kbCIw5j0GR
i6WGrTrPsfdACMEBXYlUDMe6vRlmZ+MhPGDWNo4aUrYvIbMAdshFYdu0OoibA25X0abMgKgiHfnn
VEgmAe0NqaI/o4fQjTBWcsfyFR/GXlx9DxoRigltkACaAPAGs+SPZvoNieH+rSm2q6B/I6P5LPhV
Iqla82CNqNbeW9ZN/00vcl2Sw3xp2FJKYJNVlsT7mG1C2bWXQ6NGZbCPKpmHdyjsZQcKDZ1ydjf0
s7vJCLh+Y5d6yrlsNO2HFVEGjwvdAAhxJV4A1vQW855OwB/13wQ7Es6J0aHeSzqXLkICyCwjQsgD
Yoo5YrqlPxhOLhLCsNHuakvYLbo/unJnjHPnzXlM8F7jyP2oYsvFLxoobEXvFN3GkQUrZugGE2uB
kaaBcY7Lia/RX9HyRCdHo0toSGgGnLbKm36DKOUxK4umiCnkBFPurOQht0T4OEeM23Z7Tp9/vO4T
2fwO1Vj9PvF+jTkL3uQFNa1wcbZt1/PkFiCzuklLaYyheQMdYu/pvHKGir8ypCjIkbXDx8QU0AFR
tDyOMVW9ssg0xO7J5nEYJzmLqQI2EUqgFt9hCZgk1I3zCWoqnr7ORuniI1aKXdwj71+HJQnWM94/
VCwSbNendqqOaPwyDlqz6lyIujzU/2oJOzBT43dzWk21dgWUCeaweOWLAgwcEIzTfWaimBHhDTL6
vjQiXNhF7HfeIzTpLkQuP5Yu0wh6gruR7PcTEltG6eAf2s1UoK5/eZSD80XFTC2bR5+9lCgOkbck
GQlYXO4mkULaGf8H7dfM9sigcc3zT3dDB5HMtpJLy3IfM9p9mlBaML+b5LVdGtGEDGHMEbbotUDi
/VevXCq8CvjL5qcCaY9zqLg9IqPqoeOmDFhr3kiGdT8K45QQDr+lFMWAF6DC/TMylPnIKZw5mdul
ZqcDOGK/lgtVdIN20Zz/wNENHVqpPpqEWxwXNOtix5ePqXocDB9iLJslQNfU5rSxr2+Wy6M151H4
NAru/ZY2PtpPedz/eYV8CwmWrp5gW7WDWujVazgGAIH5tmvc+DTb7mevTet49AsGVDHohw3CF/TN
RObIZ5Yw4mNk3Y8XYShvLRy1Ep5jB5oZZa9R4OjcsqyHep+P7TdMNQVE8or/ddKpf7Rhl3jWK4XB
ViJ4hFRYpxnnci9t/AuPLRTkZI6zA0tbK+AU2OxKqdImaohhfVmElMypQT8800P/V6WHb4AfoA0k
1fwW6uojcRaBdgUKFTO9cd2iC886bBHh+JOesg7nJegTp1GO4/H985fpMzdM4TztJDYzSDpiUJ26
jOKCetla2pUZcklzL5fJXkvvQMMDF1C9a0wfYcyVkOOQ1b1vPoBYBo0Z0cXp42/9G1zfM3JACaGk
54piurHd3PjedNk31xPcGoKDqRFDCyvued0nSsMI0dnCDrk8u+J0OKDwyBeEU9AaIWBIbp4/glnQ
j7cnI8pfQZterN4TA1XjRx+16Ez/zmkWnvpakS0Y4fkNh40o9J49Rh6V+Y0BEp+AvHSwWs/75lbO
tZX9HpL7tdaRdjBXh6XL6Kzt/UrPTaYz6YqAjDGBh8TLXH/PuvQ5/Bghl6VvgOzjnYwWzkh4cyD5
hBYwlBuC3Jg09k5kdyQ43grWAevfgnNZ794L5GyxyBgzVNF6xXnYcJRbSULRz17Ebbhu7oR4C0Uy
+22TT7DBTfPhuD4DnvSW49wsiVb3LYZvXGac9LmKllp7pv3qmSLUb3ZvXvY7b9b9IPLrVcLH3xFV
NyPwyFapQuNiiL1FHf/OSe49rwBJs1KyoMpt6YERkm0rlQG7MiGuP8tMl5U0sAsBebfxk7Y47A7a
AgLxLIv30oT6LwttSQuBOQlf/++Wat311FLXSoXXPoODPhrjwHFHewa0u9vMAVySVEo+yLc7rbds
fNJextP0a4vmZpLhXSYxkRlzEOzUGfvpB9KpaEwuwyHHHUgdtmKpU8A9mofuesPljjaDqFJ4ujtO
IqSXQJ6+iYyH2G+iMcm7IgR8lGotukDtTI0DOWBTxF8W0t6eFCtCgZpTrqfKhcY1xjUvqC44iWdS
p2bS0j929In8xGDZQ9yQx0Xw5fJKjBlpOWCGM0TFiIG1fmAiil4LWte7nvYigm/beIf164LmHTMT
6vkwYiFBkVWWsklNeZIVqFUsJxYyr/9PW4Q3F7EKvfvcSrATPU9Ff155sVnR5TtlINvJipowbrFG
OPf7Y2KQryIXE0fN7HSTG8LzHgFnpRavPXkpCn3T2yLP/OT2aAq+rBKTRCmsu3aFLqFmsjpP4OKA
nbNY2V8//EwiBrXFqlShQuD9H9RYl+8t5YcPYFnrm437nLPh67KH/SfFHrWVdG+fX5TSuuUhsgG7
iOhIPb2tTmkhi8PsyPIN/IpcHRBKTD2ZITh1wZs5IRHUrTA+vs76FWnVxriUKmz1mEerbZrtoMkL
HC1SsSB+U29RqSOcNAZxHq5FE0bLvUEvOlfRYGHtiZZN6rsCPoO/5W/aaVAsnvfxrmoG7UKpp0fK
YGfETCD4J65tBYqcQwt16hQsX9G+hr0RKRlszJLHGgZJYUR+XeTtt5B8HG1PUD3nhJjAPkn0TntP
iNZLV6zNmM4Qf+ML848rhhInDnYwTTmuupFv2/200mt9O1u0AE8Fs3OYpHo9AjBBHQFhxg1FoCzu
GvOan/zrHdRnFkBTJS6FIMKSbqFfudC7gfKdEiSJvI2Pu3/CsTX5UhzvS3xjqkosjfsuKBGLicyX
WsK85Wn83h/mMIA/4mW2EEEqUukVJPGOfRAc1hQWBuKmOJmWzp0BdS/q7UweCCCh9FgfzZQcmLS2
FJliSLM9TApfQ+DP1hDQmQ/FFgKDEZmOc4997VZuawpckkjHvxfV5SOWpAlNtJWG3IF9ipFVkoJ5
Fjl+8HqzZ71IgN4SdG0gnVYoh0nl9LfeaZ0XF0X4sNu5LDMIxronExoZXVXkcXq/2dPuuIVdKKMW
YDd0LG+iTbKdy6d4AFoE8M4AtJKRTiMFtmfrIsJ5UlIvwGMhNAoqSsLXTkgOXjwMd79S8qKK8WV8
cSbO7X1/QnXE5iXCV/Kgb3UCQIlF+kQEucWYKGBHMLScFEAqMAzZfevzFERt/0TkUtvNAO/r4ig1
msuZ53uCK+9FdUh+c/ZR6ZkgD0SsUTtB7VgKR/QxkqXbdWLhLIroQsVrqPC4AILjgv4U2kNagb+I
i5qIy+YNmNK06soVJsre9VT3FINr5WZmlDoK3CgVs6ahqCTxxS74VumXLPLc67Mg3i4It4Zmd40J
DMUNJ0G3qg7Orp//JkIzQ5nUcEnWQ9KHbs6/H1470kjfWPvHS3ovBZJeQxduGjaKGgdiQyMXRzQg
DvR5dErr5PqjTza1p7kfDy7vjpxMG3zgIWACO/08iqiANIuE3AKxz5D4Z4jVoxTf3+D6QL1jjrX4
VJxgaC7iQEIyGHSIAk9CV3nzk/dnB49LMHZ9ivLswZctiqXgj+hT7NVgviDXFQIf/13x6j7jaGGM
iBEOag6Ugb6FgwY+u4LxsEMEWjv8ZYVtigB0wZngK5s0oU8+AEgFEEnien1/9XB5ecGgBQk1uG64
XqrzUOOOIYmAQdaKx/zZqnNQhV8xNFc03burFt9gj9VXvyReM52ynXXpbng0KLP5V3ZJXovdIRhD
9pHsX2SJ3sgl21TMGIMN1hijrt/JzXb8+gFL+ot07itdJARRrUrWlI3vJqcwJxMXSaxH69SIL02K
kcQpvohTxvaHs3EGlldSjvRq6HZjjvk+NCBipEkjUWN6/IL/NiI7WFaqiQN0+s7UrvBnHDTdwR0z
os49gjl+OXCBYbwsZLUOA91oR6eXIIIyQ5JTU+SfrpEcJXcZhNUBLgacQ2VZuEM1eNryVfTS5u1L
nwO3fXnj0SaVXHoEFlxBLv/A4OaG2IkzZXx29dZeBAIsEwSI1D1/UqAOkG0fnjMFcvZ++1sBam8h
MCx4KM27RwVGgpqm4pOhh+hmYHZXZvc0l5s2RVt5f3difVO9bV/4dTlOte4VgsH2ekp6WXo8c4y/
KqUp/t7NKGEkalPRQlXdITg0KgrpYpv6HfZ2BsoA/edqPJET1PbsyJw33F8sLfHwcj7+5KEr5nP2
0SS0mKh4Iq64TzShZ6wvbAlRv3BgJ1JY5REV4F4oddcQO5NJHe91TmVpTdMN+9ALWIr8ZCPRw1ne
SGFmwa/f4wEyypo5gpbu+Xaz3ubCB+i51+SChxMR8lVtb4Cp+uy9Bp7qQ/WhI+5ARvRo8q0GTS0+
1PNqfH6RyF2AI/8kGPJduJGLEePR5ioYtW3y+xqySZeRhYbg1cHs/7DjTu9kU7/XfLei7O1e+Ymc
2C8avlMTrAEENllPDE1oXm1nAY3+B1VmtbZJ54omlRc8idWLygEanzhGwW7b4V3Itg9p8nBoghqw
p7Mo9xi7Xi8NfjqAZ6bsYfRzfhruirPc3n5TrlMc7q9GaRkAAAthTLA5SfSp86/Vn0oDDMhDU4k2
C9F2cuXtKJQDfNF20F5rwRYgpX4CyZvUZQgAYuTbli6kGzeSc0N7R1b14CccluNzBTOIf5lMfp3L
5yjVdyLoZGlXYEHthsD9xC2U5e1f5ICCY6L+vFivDEE2sQiiz02vrk3eldwulVXdqDr+74V9VXj1
95bwHeBbtR/PsVUOufvaPV6CoKgvx3pJzV0pKCwFvxYjGsvyixqfdILjzcNzia/3lsuehtTgEFio
JRffGfWMIKLjANU5c9M0z3Cot8ZMFJsAbSN34SQ6PX1Ugh5S0bYxpyzWcDBALG0o1MQGJxi3/oiS
p9sUT97/w4Az+t0fOrH0O90xdjqvyshhyv3EHkJIeP2uRdy4SHiW2uLL33dl8Nnoh/SmVnj//X9C
5ONaeBf+3oR0qwuSXzaZ3NqEkKvanUMhX2uPT927aoUIuhJsQopeDcNNZd2rW1fS9k499qaS+eWW
pvv1ApweN7MTCSRCBSP51QSx9s+Me7qIB64J2QqU8k2Co32mXS48VNKq+c57hXyd6uv6FU0sJdcB
mqTDSe+b7PMWa4TQCnMHnAOX6tEkxKInI6DdebmO1SmkC3/jN0hH5Glnad56tBqRpl+xBLxu75DF
FrHNXk7/dpA/RqZLiAgzAMHAuwUQSmy03Sb2DHj6BGgbJo+MBelbq13HVTQojDJvZGH96+OBVe9Z
BYOxf1HQXSx4bK1qa/PNlbRhTpOaTJb4dST3cKqvQSQZhVNRKEc87im3ZtbHh+hhWe06NbhovQwu
mvq6iganhthZzoGWZbCMq2y5kroM3G2DOzpfzdSetZxdBkeimdQVHltdnIwnT4yeoUcy4kxyB4X3
uJC/tslldiRbd90UFIY9fb4KXhKvipAxJjGwcDKZzbmGOHZEywUR9S4CnGrusMW84OZpa4FGu9+q
HMeTA2Ew6Rpj3lUTjJNREDjDFSPao2lgjxF9Qti+xKMY2Vev0a/PhDiA6RWv4XlkI5iq6/K0KM7s
7q/Jdfb2xmdZVX2S9KgozDs3sYnEtE1WiMLaadZviqyYsrhDhDcRd1wdnAApOB8bwsifIRp/L6yq
p2F5sjLYeA/Pdx1Z8OgfZUp6B/lgOlKZyHuPI/+7cwj1dE8rMJQ0OzLThGH1bQC7PmYeckL7Sxrp
j2ktmYo6OMgfXrE251AFQ+USB6pGjtdWxW2JyCYWQBcJh8R+3kvf7s7Emrqi+7i220EhJuOrnDr5
jrvEWmrINC6ogsj3pwHxhECVZ9MUbxkRBlf9I4ydob0dUpvZ49WnaUvAbw4IqIJUa4cH5S6bTh4K
+Zudtlo4ez1xe4UAIq6PenwL3ikuBcZf4s6CKTH91Izc4peExHjBxsvyck1P0PbIScPEOReHJgfs
C7c8FrYAH+eQKcZdzQmVtBf55fLYNmetr4Dc+O5F7V6M/Q1BLvLOqFBNwKMm9txfAmCA5NQUGPlg
ATDUKcu4/ygt3Z+o66/vzci4WC8e1S3HRco5M2Uk+/B1PEuiz6Zv5sYSHkCHsUEEa0hcAYr4xQI6
Q70JLiLJY83gA3HpKOyraqUOblENP3FF90zRCQGGfIHiK8xYAP0CZADkUFLYooIzww5c3upnhn+V
p33RkUYQ/JVp3rzOTETCvlC/o98di6uqid6DrLYubv7GgpUVQjXba5yz8ro0jeqSA5DFLWt6URM9
ng4QaMQYeZzkzz/npirsPvSGuXTbsmO3Ut3KsyeFG6ERwGi48eCjkgbXbTbpbCGMtnArVY57+mZg
9Ax63LzkSnrrGH/AaI3aT9PI8PsXuyVF9H1J4bZ0a6QKnPh8DqUSBbbdvc33VjTDbdo8qi2O3kB2
6YvzXjZRpBCwiJF3VXfQK6AHVC2sQqtpVGOdemT4oZV+Gq2L7lyorn2Yj8zEUvvowNY/COAhGD8r
VAMWrx4ghHTD3jqy0+GoJhK4o3m+WrIwsZvrt4erydu4A6fnFEmipTrDs0jhLc9lqx2YlhH3ZjWT
gZT/I+omXd8KoMehVl6zT92fYsX9NtHh0VtLk+c7Smx3qif+8jLfV2IRPZ1aXqJDbKJA/pZm2GVW
D+LGZBfx3QWcW5/YIRFX4h/g9Qayc3VETre61LWAauN5rCAh+1M4BSg0hiS/2lHN96LSUma31QfE
vtoXYCekFjdxPTM9lbLCaqjHF/mPeIDMY+gqF54ywYuL3TefAVFrftz3MaRbmVAYHmU3JtT1SxgN
ed+X6x8gcPdXI1slApWA0E9Ykc60z9cAPJjWNsZ2agOonBO0JA/5nKQyp7aAH6SKY8FZR1SdkrKE
65X0YF0aVtIdyR00tQIDEz55TCJm12U4OyzHHSye8HGTMYA/OUmTDFBfft2oJgM9bqiTLz08Vr3n
o5ySOlN7MRmdRLNSdCYykKqDaf9tblo5OXNQrNwpHXTAPLsY+TNNf0GjnW9R/f+fLZJ3GO8+1N1o
z894v2XsPfhNL+uEz/O0J3VcTahK21CfWgZy0m4Gax9ezgOnj7wbqSf/Y37ZVVBKNI4zddJMX5LH
b6uD/1YjupqFQysWIUbLPHaCukLbN9eQirKMHOM72gYyLy+kIzFLMEnWBv43dQfzL+HQzoXan5HR
EImYNuBZkQVF4MHSA5f0Yi0NnFSEniDvQuX+97bURKUmOgAE+3vs/JaDGZ0mpZk1QfZnH654jM/s
XntrBMWK02YAbhV9B5WEVYvqhqoc3Ev5zKruj/CZR3OiMO16A6Yb7zjazya1iFRKLoeYUW55HcPf
zPRWKzRBawseZMeo0ALWyFLjcRMABAgt2JM9x2+SWII8874JCu6OuP33prjaCQdvFfJI0XKtQ6W/
XwLYjQht/yGgf5PSXe1dnhQSNANtIhtexDEJJeUZl5zwFknnrgpOxe1n40X7ZjmYjr7APdJldqCi
BnOf0gijUUAKqe1UzSLohOi3k3eurmalKS2AeHhA2kCUhalR7dJC5c6mXEFF7zqe6Z8KGvcepCfw
kiQA5iyvWzp1qUOZtsaPFDl6/ArF+FA3wmLfe1PglbbEGb3tekNDUv79QOq31di39TigCF+n74Mv
2LM70x7OB8OYZ9xUDZOx5o8tqxeRJE3Hx0Qi4oDNWJso6ZFAaBiD7xYdms7l6Z9DIcIK4NPyY877
DfDxZxEee2r/9bcG8GtIh0mX29iBbzVLuwt1p5THFNU9m0sG/sfoSQFRGbZVJDgO12IyzyJRc2Eq
b3gXiJLONxadS798g48KGnIkOYLXPNUCHMzwcH1EbICzi/vYd055kIBGQR3wVOebhM6qtUiQmRJ0
v2AWlI+geEEvynuwpm92QT0K+1b6sZ2ahzXZ5+4lgxwPpcS7Y2rUa0K9V5SYLkyTZIcSTDrKw3pA
3V3Uc4SC7pGDTKJzuzHtu+L+jZX/PYUDfssC4s1a9iMwl9NmwJVzbdUQWC0iiBmYTQfTw6hZ0nGp
T9X6h43J6TzWp2mkqHzis6K99mxEpkV1C1Yiixb6DXJBScFOAGi7GZc+mU+r0JlPm79hQl2wWWS4
HvF/xTuKC/CxnUfvDTdNNJS0y6Gt86uxShaj5QDX3FGrD3LBNg50w+aUlRgOT9CL2dcGsuWBkb7T
bDnMWAeFQphwDdm/0I3lv1xrvvAwislLeCNaAI2RCEaCa/XaWwg6pPPZCPb37Qo+yKADBz2GTjbe
IpUMH9uCjPRIByijAB48ll8LB0qjxu9R/NWeg80ZHq0ELvr5sHqpzBsC6jQmz1jUugc6cj7YxwLY
gz6cehaZUBmW7g8fZZn08dnqmiI+XYqpVmL276IJDmXUf8UPgr5IXgqEcVEkxTAG0zzOILHZsA7t
hoqDreQtsoqki7b12pnhCZTywduBU3gJqHYGlv0FRxEbmgoiVnjVX76305s2cjlANgoaWzfYwR/J
M6oNiE5zPgbaJxtxjMVtoh1ul4UweEAO5qhWF6MCZlaC+i/dA2zv1kKtd80vuzupARW5WyA5muZm
BNoFNUw1iP9gx1lL8Zr+RG+ur8N/UbHlWL3De4gBUfVy68cCxIUOeDCO6ovUfCcRjMBF4KDKKY59
Vicx26mU1fAr1zg2ZfhV9vHZkJNsABhYx6h3PXaUNMFHoro64/dBoNibMbxpEW7UQuFrcKLCnZey
+NFoAeEy51+ZdhcsG9/eoneR+OYhcbMEdjG/inhV1zriJMlwlpgm9b4Bjhek+moRGYEfYTUdG7R3
WXxi2E4mfbKBYDpwFlmn0GTgtfYPwdSgxOUWfEUagGVWj+HULgEJjj2Vwug3wkHjYZPVjCgL8gjX
ZJmOM50vSzuT1GGI+dzAvHy6Apysrk1VQTjNMoHuMPuns3P//Q8UktXl8olb/9frIh7hPtEmFZhr
iYpDmg9EFvvgv6WJiWBfAZrEjUI1MYTj7goVIiG8Hju6FVy14xRslLjPgAGcavfDAI7SApUv96DG
g8OjHH47ZTy9DsZbo1BIJzvkRsv2n+x6t80GBm5uDT/cGGjVwRKj0qdrKAXREdAYfuzG1MoJiYoS
G3ZqF1eeAgkFNBa1B6kvByfQMWiHAWf7UhbxrN9ZPx0eJoMAdjREF1DDqrfyXMtbNu6L4Gq+iKYM
k36r7Y9tdvqYs7CKMYbPWd4+bfTsQioajO9mbUYV1MuqQEIOPdYx0ddgFqqM5mvEOypdDbBsXD6K
n+3y7sKhT16wVhwvR7GDK6qsYw42fWuMqyLfoxYSzw1PsmrRQUoKpWWwW871h7EpsaYkSACfPme9
tqw3zJO6FAx89Xf+IvK6myFH6kqoUIfrbELLIi4/F38P4UcJ25qGQAk8WQ+N7n/gcINgVuXb1Elh
O2N9wox+U5TUNY5touUh+QG+Nmhr+BdKrzZYgWnrR3/2wxrSeTm9YbHPe0MpRw3BPZs8Ho+SlvYu
zIqrpbrjHuDIvS/GyMLIB2cwAB+Zr76049MeaA7eZqm6kuUZBI9/X+4i498S8sm62vV8E/kEHct+
R9byIZtWvd0kcBwfoddalrMfUMjPmo5s2HDPtn2sHW2Ay2lD3XMwOgnIykl97PDCR7DgqoQo4W2P
S/izOioe/2bmfvuzmsZMbCVdprpgF1Uydq3gOypayKEPhQ7Lg99oasp5U2bRLFtFB8KgT4xf7m7K
/ZVcBWmb73eAIU3y/XKlmIHQYvNmE83mTHEqiD0EWh8TSeqVLLJtA5EUfyzvum5weD68t6CTgZrN
zMWpoILz0YiU75xJXwVvfZaMtpb2ZUuucPEhQwB6c2GtoQ6Nemz9w/2FHNkj7UeZ6W8pfsGRYUmc
4Zq+qBUxWfrWb3Fw1JUv7VY71Ts8pgVQdThcRFLAsn6wiXUkzCHo9yMEDDdy5j6YzhZLHen2LIHa
IyTur/Ijy1vgl2dZLLrzPhSgySy4Xm72PssYgwZlN0f4I8j0dhmZBbtL+rpK1TBoLlPibyrfps5v
cbg5JSF227hwhrnsWKBxwWVfgV4n6SGEfYdyRvHpTfePdxxF5Xaf2ZGnq1ldPB8tw3H8bAcz9f8k
VbPU09Ar0GlEbqmLogfvz18czB59JSTbIJM7bRZzAaQJQGCX0+h9RBZG7v3bSPY9wsqhVPJfU4Xv
69VcSfNNedDWCGMXezpDscb9Ij715p/oxh3ylNkmO/Il7ZkC91ChhxSE2iRVbf71LdSl5WHKs2x0
WqEhAMzDwf4JC7JOHfDGXvgoancRFbz5pSukymZYi2A6gQMOBB8ezOrvl7czlXcDxmQ6uj7nPOxl
kxgTk9rRj/vryAU1yyJxFD2rdhdlDIckM1zYVbJDVVbdjcJxPPQWjwwRbnjpxwZmTASVAt8VIPc7
qb1C9dU2G74HJPQtc3qB80JOx9UiSskAgINXVWLN30lSpyf84GZkx+7gG/sxGrHNwTG87QTAG4sf
OEbR9rfogtzFOfQLYQKxiQw/fYnZFvGk1+xH1mEM1sdrHxJ185qDIe49O/0rpBLdpeVAxYNx947G
MEPU9WHF8dsi1pM9/blYIc19xOyxeWSBna5CEz0tbgjqMVkSf04nhgaAwLYOEC5kNP07F6fE1It2
n6lpWr1HMNQOVNCrf0QDYtxaZ76zkbyAIxWfrDVmIHPjHLp1HNW5gEDEtQgyh0YrGipPCjh2lMLh
f3MdAT98st/VoFkbu2lwWx1x5+X23VJNPSMH7UXKJjrCe0O+6byVMKDu1wD5XJzhBCwse74Sg3sk
UDZj0l9JLDsYkxGw4jnXGzOnomDGGAgFb7++e/ckoEqyrtlDo2fohsgoR/5S6BA23Rju8eW1vUgU
ankNKAq9njKMUA52YsBKuTBVp6BJUO+JIIf1KGZvB4+tjpbzu5WCjnl9lDtHZEMiF5TlhY1DISli
FC8nRFrjHlMEq2NPhbgVZOgn8rPzYAQ+Tzt4jAjoHuTdD18fwh+CpPeT6S7osAX0sumeX/u0ILa2
D2PPddDB4gxFDQ5ctvfqbLgB/OYDRjUXA/lU8KIaKte7BLVjm5yYbpdM+qnHi75nFIj7YzMEWLO9
tF13d+OxI7ucvLo3/urrXOoaIxmHi3sR5Lmd2IofvtAUuo8ASlJs3J5Zo0zd0BMh4uxvbFs1lxPY
jeLgewC+ZRKXCfmYBBIyhih9UjyRqJjVVhmTV2oFWPH9jVqV9FCXs6JovzthaYXdwIN3eX/rAOTd
d3WJpiy8KZpEwqAlCI3ats+CLYXRBcE86i0o6+9ZdrnR5xmGoB6AX434YdEF98jzM88WuwmXJiEv
mPw7kP/kFIKqMEl24LnGUNOaxKFtb2+5f4XrshJGmXe7drnlu69NE1E4+RtouzphaNSWgqeATrfx
sopNSc4mCliTvrO4GApXSwBYO/Bzt5S4M7ZBRPDjPwFGGOxfgNkMs7lEHnxNIN8A7TYQvn7OmHM6
eYxm9AlKst34WqdzsbtSig0QJjnHXtrvERIyMayrh1WG/rc9Jy90anT7Ku9eRLq0AVEPna3fwDLc
As+o7R/kWwQT1VvDTFIn0OTRvygoYl3KiFnMaW9Bm/lcP/6Jx01C+zABWKVcBrlgk6vQ4celTSpa
m1+CIqG9BZNdp3lQrA9LhgqcxbZ89cXdwsANlkTX1zB1OKdcpNP8D879YFMmveYHQR6/e7pQm660
sscLo28Sja60zixLrpdUYRHoRhbI5D3/QBkUXTuDVP1hXiAJV0xHtx2Zw74z9NnWY0GjdoQbMv4v
+eBo1F5AyV+lMIIX4yHBd+JqI4fiUv2ALAVbyv4GaGHt7+JF1fg5wNTID0kZGmwe47u8f91JUtmD
xI5lQHhjHQP0L7UVg8K1speEbAcTY2ZgwFnD3k7pbkmtCFYYsUnCcZRxN8NjMmphtN/lbri44khX
o/9OH9dEklT6nj4sLfOeBU4kBxO2F+Zc/1oaEc2lIp9ddiirRiL/XAS9kUgsKcmKcEeX9iivqSO7
XlkZ2TWVrddJ6EvJ5QdXBBIFSbk5KBv4zSFO5WVQWSpEor6p3eVZbPJKys+BUycyY1Fo6MgCFkPJ
y0WEalf8vuT1s6H/jsh/DFuwLmUh4kOXx7adCof4t+OyWPn35BGMxu0o6meNEU9hALv47XetDAwD
OXTddAHh33z4ZBIxlioUXDGWhXfmFJyVOLGyqyZOHfg5TTJkjPlIRJTOhz2+db6/js7ErcB4xVan
oe/9bn9DR/Tlsp84Zlvg/pEGVRAoKaeKMW52LYN6oIgSDGtmVc4SX4D/NKrtiWPO8IikTwtQGABC
vabNiQ/0/dzLXrZUMLEwTFpK/3samiL9rBXZP5SwetSNwvagfQ5Ay6ETu1U2LZCKwJ/yHBwLUJBy
vRlpWovberBT00a3ETShI4L1RIVJx2UV79hLok3gj9mKu0pqJ0mVs9+6X9Pi3/lyqKDBKGINlwPO
P/dw9/ecV4AmanZYwjH058PWdR03PGmo+gCWJ8yZMqA11lRtW0BYR4A0dP2M2QA6gMHE4M8WZWcC
9ZBlJRB0g9CrA589mbkFQV+/sU//hpNB+vSLfgxVIXu8ROYRyFGxAcajVHPFibFlT4ohJ/GJYndT
PhFuVyMm1X9dj5JE/UOgjp3Ab4Xb98krV4HLpSvGJ7j3Nbn19JGj27WpnBf1NSKuihpjde6LQpKs
TYBMF7h/JP+PRVx0cnfKyNrXDd2FtGLRtE1f+EC51QF+F3ODgIxj/rGhrLwTpvKN/Vzdx28d6jW+
M8KipKimOH8JwHtRda+zn+26CjISC/9NETiU7REch7alxI+6/MAToFn5Sq6txhDH27nK+5zdDbK8
9uiFKjmswmTUB9c6qwullRlcoR6Ajdas44BPkk6jADVVnY0DclSCrEIfPYAKTYTcSIvfxRTNahGc
fyKnBodoxZvDgGZDeygV62Lm3lAHjzJMIoi9nKqHmdLKLIZ0lkMqZKoHiXPWTFg7cpR8BB9qI6X9
DqjhvQf/ZbMn+0a9mKyEPSlgYnvTyW/meRfwBjpdjLVpvvWkGOD8jwGuQgO5TPueE4e9Dpe60EnI
HF+tjyR9ZZJE1DBPFr5+d+Yp4dqkRkKwpM/te5ngMAYD+rGOmOqjU6zQ+/wi994c1ioe7NqAb8O3
dG4hSfd+6tSulECoZjK49hE8hy9bX/xIL895tsnkwv6n1S3BQv41pmAsM/DoQf1JUllnKS+Nu8Px
4SlqUPtDJeJ36DOC/C9/rXUHBVhD/hy47T3pBjtCTmTIvOcxJAf4vNpCHwRhTIRZA+NxLEhNB9JQ
BYC7LGfDOk06abv2GshHWxguSCKTLX82QRI4Rr15CiU4tVbA3UCbit/vxHzlsUPM6Fw1OpYnxlvy
puDzy2OdemZeVdZIkdJA/d4SUsC4ziHZX1Gxiou6TcL/jgUrxzPIpXnCqsnOLqb/3XVHoITInFgX
9bUEy2dT773HX27J98tkVqT5X/sAZZZNhs2iX+/2yOvAK19L2qp37bsIROJtPm2ZLwrZGyousULH
f6qYstv78nRceWLxbEqp1RqwzGkW/DolYEtbNco7Htx+tLalp1E51HZZlC1KJot4YmsDs+Ts2DjK
F520Jn+rnCxX/ej6A/uWcrqwANg2sqlWkXSRiUPtr/Cb0jCDtLMrnUbiGqllHrI9cYTwoRei5/h7
aA44X1xzmAvQrMtiLlKXIgTFK4b2nE1ISHPs8udWUUfTZ/qHI89ejwKSSiZwXbrRBGdI+Cefv/bq
Hk1vB6U6cHtE+511yGjfjirV72SMOCnWx3ALJsIiPnU+ybM/iAfJp3uRGTDmqZ42Xncz6JeFBMjP
AIspXJtx6YxP2TwKccxiOnyQDwKH7rZdZALD4iEzxxSIpMaV8kgWOxV8+sp9MmlVQRIR0u3pnT9g
RO0WSExPB3qJpMtWMnmFqU2SwrSTrGxWJPCBjzDtP7ZfKcdDnD7JZl0j+0sope3nGBAy0p4Pw2zM
qVx2UKiLKJZkz3RYYi2yu7faI0Q/35qfL8ji6Yi7qFVsJMgbnhQ0y673K7ZEWaMBr0VL88mtj1HZ
dKWFVJz8cQ49L0AjR0SDLGVNYItBae6ClHjypRXnzegL1LW25avGqMCt3HpdEzhkEOUv/A9AAUyV
D+pwxiOlSkxaw2j8bqykSxP36SPj8fAH/nV7jIllyshZEodaU+bXv2Q8Wtse56VwhQcma9Dvpssv
41O7K2NaCuL9DEeUpXJn9F6DUnJfRyS3GF2FSsbz+FKH+rD9q/dYmFrSr9TmfW2mEhvwJsmt6LL0
OuVTrf/9I1869BuP4ZmUYlkHB05xunfKdbEphTt7c1ILix/RHKUOvgTY6OceM6gVMK6Vl/jSqwaj
a5R3sxx1nnB0rsjbHmS/cxnJw9BiLPGPGLTYb0+8wbTt+TdjlZrzJb21G/yizD8QXwDhbLDpc44L
8b8/zjA2uud3dn5GZNqO/cKa8kc1wz0Y0rUE0eKQyqUN3XXSM+p0Mpc+tX3iO0qEXkcV+O26KqtK
f++kiq+n78tHY2QENmJ0eE6iu88xSJj82YHwT5rtbcnonc8WW0XcpzMbbBckorvyZzH28g5nxh1h
Z0WXSYCHf19ZTPSKi/E/d5J5xfsRSAm1L/r74RLVS5JxJc34FgrhMX056gQLtStimPMpyVusNsRu
W1XUk5ZCzPkgZK0V+MU1cMmdtE5JUJ+iVVYSdTtXopQ66pAGt2l043+GtOFcWPoONB1UHnVFoNMx
feIwMJfgo14ZuOy3wppcCgDmEJgSfWrjt9nU9IZdmoHLGeplo8YThSTmCgn4+q6QPzLinOa4F9e8
Ph6Rpz5rCoChiBWoV8HRo0UodFAgXnkHdc5KvRzlXkh9wUbcn5SglbXAVxh7b3BnkGfJJpFL86Y8
Tiz63qpwxgWvqp305PLR19fifkaaVaQiu7GGGNoZO9w/sFuDcbrDPGernaSNGF8bg/CEY+ybGFJB
D7aF/pIAOcVf0eUvFvzaQ0DO/jK5puFbYMq4CSspTSnZLqA/JiSPVtZnjzMrNkA6foeGd4sWktUR
UX/cR2xzEqT+01eS3fbPUgdNVdEkL3s4EeGv+E2BZRah26uOOxbL70S1wBPb9KzdtwXa+5LYkkNu
9PNrUs32aAR6DOE0vdJ3IphvonzuLL0vy+UdB8reSpeyYHaxJGCyoy59tewk6K6v67Iofo6wqiOh
G54GfPqXtq/lG4t2hBoIN56DwLfhQJm24tu33EOL5BnNLfM05LvEJE90c+F4CPwigySKSMwlJJFd
4N2FqU5IOZbX4hn6n77dP/fKdWAmTkCyWcsSnRs7qAb5G3H5+wIrcMusWFca0xD19rtKcrQVCxNS
/9Pxonzw8O/Yi00APpW36+mEeER+tk4vZziFiL17L6pE4p3ofB6bze4iBEBtyQ3Nq527PYPAz6QL
6Ons8l0RyJmYfeJtQSKAwVTjzfKMH9E1lNbkoDWXYjcjLZIT1N+7grzQVMx8HctJcx6MgFt+0oyk
9i+Mvrx1LvxfEJeCkmtJtK8rn/J4E4OD2AgSmyvpvXJHIJ7OD1dzWceHIpeFrpAWQYi5/CqOGQpM
fJGDkcFr0o9cIYS/trl7YzL8pM15q67uZbJ6V67TrIP7Tjw/WTKJIloX0Kfl9S8XKMyIMwmckQ/A
w25HjOIg3DOA5GPR1WgBXgmcN0NRl9Z+UXVX7andhmiNW4T3EFNSZSuos539+gqr84iXVakn1+zs
GPhHD/tkdhizIA6Ocg7bi81XqGaKWRXYxKvMGwhHsov2k5hbI14MKnDIjpyDUKiD2oy11B9n4kLD
Ueq2Q9Q1syeMBl/8kI4BVPJI4TDR349Wpub4yOsHkJpCQry9IWug9JMx2llehwiSbe2BRbuhQ8Bz
bbWHaZXXHsIo6pEDW4fPvHgJ2t8PVqvxg6OMMopJ9JFLuie+Y4CSmQ8rqN+iqDqzZrAw5naKoyty
M/QNiW7L80UlaGTFlpuYbrew9an9Mu3p+O/lE7RaV5N0kHVxsRM9Wvr3ofhb0NTDyygkbpnPu4Br
LKBCnN5CNZc14Ego6VTJgktBIAVtJwMrXvnnWRIJD4zYDHri5vaYGnLBxWNAKtOuCwINQWhm/SOf
f4I9/pkI3KfVd3BcqYHCZWRuYz9IN4T+zBfVDbUJcV6r/jlQnqh2Xbq1NIBsl3ECtvPLFK/blxHF
g6nAUcYTwvEjt8WNRSequwEvNpxeblBuNJ/ghweVfITmsNNqALX+XDX011oNe+ELd7ndMnY2KR9H
dKsDftK5/AfhpwXu8PurMuX2LZNitHasSpyVtc1w4lQXmpoKP2TSEwr/BJ2WDcCkDXLx/xh5NNmz
JIQNq2sKKkcFKJHnMsdZXE0Z+hWWfpWDw+AHbxAih//vDe2rWa3Z3KG820i62KR+T6Sh+mE5wpIR
bHAAdt45YWpHEoi5RchF2wsc9dbZmS7u4gaws07PyHvX+Ip9bGAjkZ9ZuR/TSxyP1S/AzjrPzXIt
Zuv659XB+r9pWTYfFrd25WRPOUrqMkVYqnrW2PngVZhzfOXm8Y/TNVoUEGxmTv3k8b/hL1LKoht3
GOV1e6FCIKc4qiycSWJ8oumF+4K0CWGmaITG0dSTQcYhp2yN5M5XDpEBF7nwpLybcCtts5DNhbTm
z6SgwjzEHykEay+Hhv1pSn86F+r5/Rr7nEbMyeoJY+zjUCWBH2wP13IpIgqQN5Lx8Xr7ivsR7G7p
fhKWYLwfnwu2kxuY5w1usD8K1FLo4QTYn0h9odjNm4cCXiLB9u5BIVFy76+1OcmMm6XL+eWdjTiE
aCWuLK0UN10rBykFrbX1y+NrrYt8V72kH2wGDiFlUJvsXHqDuaIkNEdBtVQPiauwcYhqPLItni91
Rl19EG4UK/bweF3GiG0Lgdz5V2pBRK9m83y769uKy5GGjqhQa02pYAOqax6c7AvNFOYu5rtK0NC9
81OQGfoYrvKh2MESQopa9JvU6RlO3soSGaxozkmawaejkitXweWXFVGfcyo2QK7LX/GYhPXQH3xw
Omdzg1KGe2P1Nnwq9RKgkxLXVQ9RvqchB70b/vygu9E+a/Qo5TFAVC9mfu4Ntx2K40wktGq1S6+K
wtTCkHASqdKVP5tOpWygJr8U2eSKGevj0sTBH+/jDgmzbP6/fiMVQtfCO+FqyCHCXcHCwSmfX3jh
CBphGpUwTJrGdI9ndtDizc/T58DIDI8Mrv/dgPTqaq/y40CxJhWmpiT5LHC+ur7umz/HFFT1NhlM
AQBuNsnOVEPWM2Pu9xNNhwiPXTziJOcDjH65LMDenVAd2CcM8N1rAAjqDZz7atLtLGZ7YbGNH3oK
PH1+FMdF/LQ6IihhdazEKpMD3uJKZ6zpJ6+loFMX2TFlT3fzMpYZgAEnUkmdMercH6mOibE+DAu1
oQ7fl59j0GLh1Zg/GcMX+snXz3mW8NLnEeG+Jb29M8J4Jr99x+BtxDkjEC4NNoBPPT9kA3AnD+ED
f/PolpiRnAKl2soXSDsle2YV6jivaeWEpL4lhEa+m9u9btHPU3MWBpA5OMLDrkeQUy8COa6uKvsc
2/ff2CgSQrsTGtom3gUZoYyrY02F2A/NUIpKgyOp78jGsqCNDRstvCwk69wPJKorZFUI/izEoNEw
uOQ6iDHhN60myaD9qu34ZjJW2l1cSSjQUcAIaFNW7d7XY7Zg4dgWQzMR67ttU/wGqqO79yruoJha
SOA4INnk8yLOBSk18+IyThamw07QHn3xuhcofhIGGIvq2qjT4hAss+akhKy89LAZh4aUOkLqKe6G
BU9m9+cywSjRdtZViinnEWWBkBiPlu0ooRBLJaeYjGQA/r5eLFEzzJAJaTCMOdJWXMcp0vTtGKUe
1bRxU2iT0LLdHW3hOwt1Dq3PlZTn9qmCwKHrNyBxChX5wHA2FkDyJTevqi9sw2UDv1xmlJFYNVdp
ZqYoiGd4u38Fg7X3gQZi0AXyNRnp34wDDjqMhQJpZO8s0rKVVKIxIKyuWeORfLYccl0fVEobiKDP
l20HtF8oGE3DvoSdDPx6LiOj2Jfs/4nokOk0sE1oAzT2zzGxhAcTFtIW3mdAuhjAfU5JqtXdcxlY
TJGOIpMWYBEHPUwH1ozVnBC7V4EbB148sgY2TQRcTnS80ObQ/TVt3cm2fX9ABSOOZJgolKtsxCPY
sWgqUagzJSAyu3p1Mj57YIfEUYrsZzDXkk+NsXK4ZUg+L0ZnOpWfVHQ6ftopzc/y0A6HZm602r3K
loy/Lfu+AjsOwv3S/QD/X5fdxZSrzB1N9Uu+qqAVAniDuwljTu8eEwYO9wmKoj4YzLUK1y0tZw1x
4NWYaPfpqhDwg7tZXayxEO4EDhayBZ8ZmQwIVSurpBaBYp1WM5uIo18XRBMSQz5EqmmY33AtLalS
7PWyuaiferhIowzqtdFmy0PeYgDpJ5Q0GC3K2PQ9womAwd+BpU8TXOJuTtkrvYzRWmKQhc0Blvey
ybiHNPOkQ5njdXEOk8+kNWsAIKZs+fAfWqeo2o6Mn3r2aA8Kr1Zrftv/lufg43kszrf3BaulZOSK
NnJKeowhrc8uHqoOU+Re/JmfGBXl7A9OqvB0x4R/Liy0pGYQvbIJXbFk5xm1w3yQvpOE1HyAhhk0
2c1ZDbwJ11Xa9DrOwAafLdDnkDTuhh7J0yw2d7OtKHVb9wYjzaftdeQl3E86FYrOoV1Cp8WPaG3Z
DqO7qeduxaaM+30VbkR/LXkVPTxE1q9vnFuPCZixRLFw3FY8zFbdPz45XQB+jl8jfzfWdnIqnSax
SOqnCv1eonq7/ruOYOi26iJNtEJJVV43kBKawjU9lUu5Wd7LQNWpRPU3QAqJbLWj2ZsbbOJPcm99
CIW2oGUWKiDwT8rwCJxO2MwhOrHxqFhYGGr8YUiSzyku8baWNXesT8u4gFnUtFY32uaL4L5AHjHs
XVWkYFEsz8JcAqBbV2sdBbc1+cBc1Y0nXn0tRaE7na7XTsPyyVwi+8Z2GnVo6Pb+W2SIjHbMvp3F
5Q8F7gB6WGv2yS7MJreLVcX4C2dC75c63OEiNZ2LRlMyiyFKpi0LBXsv7ivBXJLG10uMp0cBtOjP
vht8VGfPyEzJ1b+Z9rWeHYpbtSqEG8xrWxLf0j+daw2BQVWby+s/qGJ49aTrfypumL3z/SIxvgHg
XXbim4t/UXRBl+XhXcOGjV93nooy+noIeQsW5Xpdiahcomzymx1SShUSErqXoSarz+X1lD+MmWt1
UHkcFzWYv+bVnHa9CYFj0bZjLZKuNFXOq2yuwFMiJaO84OjfRMV9qRvHdgTt66vDQZ2iqQZc13yb
cFD7UVLsc+VlscmYv2+yOmUkazr0RVEXUjb7jSyDv2nlkA67oGq6FV9VRVUrhW+LQwgd65aeRTO1
ljFXNcc+vCv6qfsqQmpL514LxXhC1ciZKd7WHzpFBH7RmJTaXQ2Fv/OZqnJq3mMF1t/dt8ObktRW
l2qC39Q3VFZWAOUp+YFMQvqDlWFQKYLnZoGWZnpuBqwMPBlTZqcsxbRP8esXVb+1HgMoDT3ZfiRP
h22EunKWBM3mqHBr2+3929aImiSst/AhDkfU4O8HWw/QrSDuGnTV6UNW1mfchPPKqu8Mb+1BWChM
efFKoZUUuJYbclB8y/1dsyyP0k5O5NNxHB6/l5n8lgDGVYAUZv6cja0BCIpJV8dHGXuKgLQBA+Fn
FMiZBd0jsDguJirBdaQ0ripBoUh3gPasq5ldXpeHLWUD8PnLhOSAVksYCZXiHOFye/oWQSmsHrjY
5xEvJ389WaqpsdNHDR1SNsETr5qMZQL1QKL8OtVR021YOPxw90yAzGMcsjEqwc10ybbz8+DFtZPV
wYggSIgnOP97GnWO7dgCLqG85dsLToIL6Zpg59COr6fvJYb7ckXq/jl+ezvi/d0vZTj44+1Bc6JK
hrgAbVF79NkmUbjCFcC/e8xW/h+8o4he50kGY3R1iTrmnQNY9pN2LXLf8l+QiYa6qKQr1prppgsh
pje186TO8eLBpxVnK8dvzg/C76N+FXYX7Uzrvc1nHe1pihYKVbBMCcO8xlK7aZEDLbwVedV+zPAk
ZxX5aq7TCGO8npxqsF60APORTfH77LpfnU/5Rmm+eekzBIvAeif50yOitvyV21RxeOlRbVqgRFj1
rQ68Tj/V0kLLSSesO1fD7Mx/Ceg1au9/xWczGETB0h15LKaH9nFd/CPDwEbZ11E79H0Atz6PZll3
EX+ekQJDwqJXDPHQkUBhvdD7wkoypmId0nVaaULqkuvul5JV42TNVu0IqsRMQCqhVNbJbXRec38R
UtNqxNYR4xzVEZ6/06hwG91udt26KK1nhFZFz9pfJ1/NdbN4ZAMjZs5OqALzw31y/W8tfjqWhkdo
EYSL8ir6RyruMfZuO2hDC7OHyYOY8T1wqxOjlvq/pOmwGF9pXjqhftzsuNRZGcTS5e0/h0201C+Q
1YSnoxHVx9MEaEunlSBNtCQSSru9GSzn+euEpDwgFLu3DRnRaKBZar/To/sv307jCHEfWp6CZmrz
JIc17Qfv9OmvqpDlu7rxMVpo8fY929Cg/u7qi08g9SFqKO3stMygtEOIXT39c7Hq459Pmc7fCCMA
lHIbSqARMJyuQmYnBt+Ahe1u6Hc0hvzsO+cFANGacBzhSZw0f05WHAfmR3apLV688vpbAELTvjim
UMKjHFWA1pqJgmizJzVFZrwF9nlWBj4qQIVWjmyIDji3GBKPh5tKXNTjFswLehObtH5ayuJ2UUqn
0zjAgz3HzlQoa908jWFfdIim4FpCDn1HJklzDeSLeYSAwWFbN1R8pI1X6r4TLAhXtmXnWxzYdw2w
H3QBVf9RmDnDqD+VT0r7h5oo8AK+yIrCTtw3V+Iyx7UwwKT76nE1C/d4A7BXQnMOx+Mp+DHOTBa8
0vdxmSulVCy5GcznKrqrMDNTBJ2qODNnDB/tZ9WH7K79KniE1mivktr9FrcSXtA3LMwvHHFgzsaD
Outpl0XmIiVI5AT2H0jhjttGznQy+NkC29YEu5o9OtcdDk/OTI4jNoHJ71iATpyfDfgKG3NB/Dds
7rMs5fegzjE72Cd5zWBpkpUugwDSo750tOaeacUVmJufCZwvYMWGu8bE73x8s7WOp/daAPFvgh8i
nnqZnWRUAR0si8RGKBi3dGA02m6nmKUgN9Zo2Bq1RnCpfFXGY0zho+VidNqFiyV/v4XFZQHVA9KY
Clc2pbqCKh50L14S/y+3uzm3ILWaSzAkowJrZoaZa3tArnUXN7niukZ8lS1RA0X1zDvycJqSHcs7
rMmMbirreVEbLvGKgiOP4uMg2F9+sAu2zDnhVkBj6TTG9Eq8ih/t77MhcH4mN2gTXd20TAhOfHhp
Ib5PnFTa1YkiLCCaEw7AxLRUzpKacFji3hdkZPftuXpMMluuHndtYR8c2vNRuCZmV5NtdWRrzbI6
4V7dff606vRweMNNkYAMoYT+9FceymNvPszhoNI9TCLCLg4chXM0KYu4IMe1F6p9mtqkepaKQfVa
eC9rgjFaPsqoOzT6oPiDFJ7RYngzHXJygjLJEwww/73S/DGpCtwLZhyx50M6KLaiV2/uoJhxiwbi
9cKxBBXLlVz0vn9AzC2aePEcvxkxf6JVZTQT8U+ab2aI4iTCfhQNkT1vsFuUuh6PlSvcHZIg/04G
8xcApFK8JZypE2sc/C1mzwQM0UFtPOqNrlMZAM0fKDy/flxPakEQOz9bb3HC+kf2v4M+EPP51mym
n3joyUbvdgkQ/8FbeWmkRLQzLCmBUIhvV0oLu4OFh+ffNZynuL7JRUnw2X1Q6TQA9v6negcgej5k
9TLJaGM7ZTy1qmtMBqrlYXBbvxOpf6gddLTHotT4nOFh+2cf3qKU7REyPYoLiLHkcWQ4v1B8Y1zL
V/G5Wy1GHq/WPoFx/zT6imnSjdag4h2ueFX/nxbWwmexUzkn87K24+fc09+x+K6ZA4aJcYLMjovf
BktOaLE6UCKHtEzNkEMwAQIXDDjUtQ96lCHw/ZglsPZeeLrJouGzNWxEdUFjjMY0UXTrLEjHGdV8
/jNwHMFCAixAj+j1JV20VjO2r5LkJd7mPr9+0SrG3qtMyYHhTYiaatzNnP7XMtxR3EvV6mKlagNX
EpNLbLz/Qk0E1pf66RsrNWHxTQdixGxhwFd3UI+PoSBehsuyV/hMhPaaks9r3knpl3U/IvrTFp0M
QQ+/XMqYr4G/qENri4x1PU6RTzvnPxozf98OhdtfQ6yZgnVaUX73uJC9KXMwbei1GxfauDStvY8G
zMhKkpmgq29cgtAMSRUd33yy29rpLz0PBYVI8YHAxjHvnG3w8qNQxrBL3i1Yx+NPRZwp0qYDfRAV
7I/l40mWYsS8yGd6O04r+7FsMQ190zZPG2zv6NKgW8znIvfSVOyfcogoKeX/pnHs4eOacOg30ozD
pHDq/cbbABVehqcFGa2/mZxLwGGIdWpey2fDCvAkTbPTZa+Ob3U4rx/0LUCJTtepkbdSmz708sm0
Xg7bjJVXVRgQqvpa0k8MQb7Ak9caoM+zwpRKBbbU1Ev1imr49lToIr2eDFdg/F2wLpqm+TfJraBn
oJG4NZmvcEEWHbOF6yCgbIMvwxtdavKt4tYWjvC1R5uibTbbegBWHOAORG+Ur5Ce0irM10kwWTbC
kHYRwxhnWlV0qzeM6djY0vZG8l7xtibu7zkxX+UQyV5GaW+l3RnXXwk2cGHxHSpBicICArIVKTGI
39WGB0N6vuoP1ENC4+xD2vuy+B1Js76gi/HngNR2iqeOczv0XOnKeMmHDkUU/E7/OJLWp/pMRENV
x9RwNoa5FFnluKZy6+T8+zZ8XYXHxqTW477LzwM8H37N/selOjzsFk2XWuL6sTcfDI64A5gMt2Dd
VnkVbEM641IBN1GSPx0dV3GrOg7tiUhaYJVEQMbDqpITK7fy1pvSPX6zHvwqUdz+aTYiu4Yw5C1o
/ba2JYzIz4BUCVyJ4WOBiGBtU/NvGekQNKY9kH0QuJG6Pz3E4fcHsNaEa1rkH+Gjm3ov/WNIaPVA
LxcKnRQQOnsWtVNdflYTrFE97UVNK/SV4BiKGB4cQHDKeZH9Y196BHve0Zhf7Q2TobUeM+BTccn8
V501fKK9MHlQVrr+YmvadUYCLFEMlEbKCqVKTAVEA7hcnkCulv4m+em7O6/qxm4Dd3gt8SDq9Rpl
xUkMfSljB7EQoJcCC6yBS2x+CBJ6cu8DkyaPDE9qm1iCr/7/gCv4Set3NvKKKPVdCeJjGi71JDtO
BMe9b53WzUhQFTJ7XaKsAPb3oOabMHZMU88DQgBoA44WiHewpdtHzieHENUUZPuAeCocETyAix6J
wrfAioER0IY+CK01dANie6dk8uVj0O0lNw3baaKxAki64zt0olFa0rjqoIyytCoBMZcMORTxBxvX
gU6Ij3p2rqhudzFjcxVS4ZdrjyLcUBVeb1JYk6lBc7hZGi5RCsXB+CfycXCTfSF1EXwZVDuWU9j2
0l/T+xAGQx+lXMzSfH8+Z2yEtt8RhkP3c1xiHFsMYtI38odM6aO9der8PVeDU5aNqxV1ifWbYkgH
SqG07nHYEka/S+eXJyV6RCV57RVioQXV7gpaPHA0utAz+p6sCjj4kD1YKEQEt2R7LL622P9IuXMq
3fZSj/MVzfW3zeksafNWipQHGZqxUu6J2byRfaM/BXvRo7R7NlWF4dziE3JPBAYC5i1OfxeafmGn
TnaypxCdnG3fxXa6k3bqYMCDtV1nE6vapi4zQcRh/3fsHgAoMHmKcYfn8qxFPuF4AzAw0WmIDM0c
8BVqX0VhcWk8FCe5eTNPwiTrMLZqSHvK4UZcFUhaE/el7ety4Zj3tSj/u3jjqnI0egyl14HND59I
zxW2p4zhOEK7d3QI8kW0KPEz5OBknA416Kbtw86a2OrR8xotJw+BU1+wXyql3ljIk+uEfanWhPOz
+djxoSQFCHmRvzjzziwU+b5RDzVh7lYzDs/k6Idhl5P5XNFgjKDYnEe/Bgd1V4W+lv4SwaD9Xa0U
pF9iqNAKKe5hUd2ueQl6rqvWe6zMsOafCr4XOluQqyczi3Qm4EaG0SI+WseEVStgK3/LTr3RJydi
eeo3fkGFO/hSe22upojfc5Rjam3fi22yGtZjwBP7it+FtwT23EnFHBC72zKzWGmd9SP9gPSLDup+
tJHUzuieaB9w/F6ygSp7jAwnP1coCd9C+n8cG85Dy+jGS7WDcw1gCtdKXM+Jmz0zDCIHn9OdoRRj
LO7LZCRKOM6pu6agAFdIzVsB6DbPSIEKXbD1CSC9HX2oHFTs2YyBu3wt3mbpOTdmKvcwwGQZsdAl
XafJ9pOAcgVAR9r6gnJoobxnb68nrRZxaqRdLTBxI1I2pvEuq8BCRmsJcRmBuilxOaG4tHBJcq5U
BhtzAyYQgQbExYz5qkzgUev89KWq8RlA2rjzlZVh9F8nH1+jzpvdkMMFvqd6G3sFyrfiyZqEehQD
UkvmSGun9YLiehhHACa4G0COorJsv9n6MSgvuBccMmvNFC3X758QJjZwnwRyehUskPYFkDaO/lns
hpCrp2iFW5T5HOWtUGlqlMcIqB+4XQXaskNl90NsA5u4GhinYibqElQySOMG8cN0k5q3p5ylMTLa
eQlvs17BIfQ3AzuI4wq74lq4c0AmI9UGtM0fGNy0RO9IWAfhMHBAF9B9/t7zyO7UcUd0SvW6OPB2
qKKf6E8MeQJLpMQ2hL8Du4K+9VjbhSmnWkqjGdq7Ik15LDrq76wQBSfYRp0QSNE+BpwZ3TR92G9+
qoFjiNUuJsCevX9OUchoarGhn48PeG6mKdiuuNmO/+zkola7aef3K3yxVUUbH5A7TqIoC9Grv5PK
JiP7E7XQcm6nKgpy0vFXBz/0U9nbttfZFnQszXbPYauD6yfwADgnQBzA/XriHrCr0qmiLBf6w3uQ
n9YigCtw7h5vff4XsmoVDsXy4dLo08j0WBYm8Fc/6N6wSQEoH2MoNGpgSccKopWGGTLAyCpWSJM2
FAV6dRPTcIu3/fLq2BoMT7zUDXSyuu/nL02StQIaKUawUykgD+k9eu4BxE4rrPRGbEgwv0mKzoZI
aa99BatvJMgisRWgTpBAt8H8AixNs6a3zuWHWES/WK1IKPFOAVvGlZhoGkuFGvW+04gfumUWnh3x
6D15sQhA9qw3SyxVlPzeMFzPc3cvDopAwIWT/QRlcMjl1DstJJPbX9lyfUqniRzCQbUpZtb6fFMg
/yh2TiHCLVgRuGBcxaBKMMkeFA0nSQ6gojHIUzdc2r4lop6XOFeGJHI6YsEBYqToJTbqKQFftT2B
ORVWJ9zEwJzP9BXFsOjj5HighTPIsF15bg9iDGE6aIFHt3pvIGmK1b//9LWt47A5v0MwjKuCuvxc
4HCj04exTJKfkva37skEWDvCZRLW+8uRyWPn6yWpCNIEhEfIsPBbQAwlgH7TLNYxPpEifYlaE32B
2iQQa0+oDg8K07H+JzNNOyd/kDtC5Fh/81Sc8idDUYHGOZ6utYioRLkfqyGwXVQrobsCx+RpmqEt
I78HnlsVTXzswQWCdcfOe7M63UkSa5ilI3uhh48dhZhG+xW0vHGsNfR+jtPWLKqy6z0NZuPW9uVW
5Nb+69uuQ5dO7rCACxRGt0K6hiCDpi/gD1c4XilfEppGrJSM7mVWbZTOSbwqRfIP3S8Tonpl4zRE
87gHlyOHvBLua2nW9nkeHDjXXJukvhr3cONcZqHWsgHnPaP/e5WnG8jaMdr09qCPZaKR2eb/+ho4
mv8889nq5gf1HayW6kowzzHZ5f/VMzH4+DlgeoAp0RKQmDGKLqaHyrp4sYotz0pdEgPs/90GnUHj
jRsf5YbvqaHgkST/oga9bNAGND5OHbhA2NOCgwt2jJ1JYHJkMtfGlflyNgeuP+1vvM5UakQKPH7G
ID+rmXqCE90WIzNyMGEfXjpLrQw/0zGuXPRyGWltMnjmOpzqrTJD8Y992vTdXj9AEOJTqDkgCtBt
YG3VxSlTCpzYy1Ddrwd0EKm26LqZWZuolDTNdp95T2VJg1dCk5bG1SSuXaMEPdedW+2Y7OdoDrBv
IWWqnJTv+fgaMlHSi5fw9urQuQHQnYCgNc7OTI0eEsf0HAgWjkgf2p1pTQybiW6BsqOURo80TDay
HwDsBJ8kR3y9FWYWCC3+fCqQfeywxlqGJbFxkL3CqNeJqfjtPocUnrGKuGlxq5y3cq4VsnfpMYjP
XC4FlIVk9TD0zRWOmn/qBGmJH+xs4U4zFdDy4Fgx5hA0YKFxJiPPd157hDYBMdnwdv7TGX2JoJjW
vLFqZ6wWOmbKFHBZSBHiM6aan6dgYOPJb6+0NArcfpOOpzbffPSNvY+z7e0ZvG3JNwkByrTO9QrC
3f4K53h3gbgbCc8NRILDDSECo/9o1SOaTBnnu00/GxZMApT9v0c9s4vkVfq+gCErtwAmFy5XzEGf
zuAd0UFkxY2kjzFih1IdozBlyTST7cuqT4h9f/uJa2+1Pe8vXiHct4afkwa3Z9mHEGd1FgINHF1s
PLZJExR1wgkwAEmAIknwYbSL3xThghvekgYaFOy2TZzAjEqLegAclk7kB9F4Johis1IIaAY28YMQ
sq8JE1zoBstarhYwa/X1TmH8gZXmwY90Bp2iYuN5RNlm1NEpmmkBdRNdgux93w0WHQv+LBRTS7X3
ov4fpZG7dcSePqwMo0LaJoazs2ZSYHJ17UXht6E2C0sFO1/pSbgZ+B3ZRxaBnQirt7S4uZCj5Z50
zPB996QyCBjlLiAOAesyDltK9g15bAbkalTCFBKVkH7h4rTk5h8XCbzBeaqQ5tK53MSwojRUz1g/
kAE5EQju4DIuWGhBh/x8236bcNfrBgK8kEf0LQ2n3247ft7v/CsJ2nf2BGEYSDBtoEsNpJP70311
5kniIIAIo/92LtCf8TMnsDs4wDeabLBOVKOlQSB6BbvbzvRhdNg0OvWBDodBNm5QaaBUTelOCIA+
THA72Sd6hk/WK7jp+joDYRNfH1UBxOFHgcbLRj4aOg0PEyM84oK+GnLTb4VZQOXqzK/gfc35V9OX
2AljB68id5hczREb9QooNDQmYd97tjmL7fIuXDAwji/syCCDPMwAEy/owK73dMNSrq/YTNvSfL3l
mONLsVWNRNeIUcVcNfFqiopwalRDAT6aekFpmGmYVN7jPpps+a2f/6hNp5FD6zaPFhdmSWHTzF6v
hfUrkjx3IEqWMhi/A8kWBRwbZG+PCZJPptJbNxUI+MiQQezHNeMOi19J0AbKeoKuvDOI6m8BSagT
9pDPQTSLmMidsG1u7jea6Xk0/vk7u9LgysT7cSjSwMyg+GSPwCTgqLqQKcsD8b08B3ZnVg/+RJcd
go7Tvj7kXS2S9q+ii7q99/c3Z2R11LDMaATi8lazflQInNEv2KD91qZ/o5yRdXB8ZvDH4AE4X35W
i408J9ZHV8vcS7HEL+DYppIEkDuwAdQ3j7q4Fv70s8FxZQQhpiQgPdQIUX2ZD9IzRsEZOdy9nxdc
1pKrO4UlTzu9O1EKCoRGSNalGeiVVuS2o3zHxG5utos8TvPUu+ieFKxrNGvbySEMkpA+8LAXE8i5
9isxmbKIPAwJUwlW1BgG6h2v3tkvmMfrahN4ahrZwgX+AWWg7Q5ihLf4JSuSJKrehu0KS3VUwHIJ
m6IVdHgLAvbmJKn6QwzEBzXxCMPhnb8xv2JNYsBGNU9XoJ4hQukRauk3bph5GDJVU5/jFwc3Hc+u
91BxitzR33WaPZdXBYhlI1/DVRU4emYDZ6PuZGRL7Py8ONtT8x9U7O5c9oyaqemdIOJy0dyAYyob
F0y+XIPKMtPwxywYfzDabShJWzTGcWCBIi5NsPkByCgJRorVuuwkje8Krz4Hz5gtT5LA2ib1iOyH
xOisxx5DSLarwFw+9imHADbEkX2b8fhgdKkC7RTe4N5sZK9XGkOfqeKafC8hqeffP8XqUwpVNys1
1W7KwxfBcCIIG7fhAGo8K8fo9dWXjE/VaFtO19xxYAqOSyaNpTnJM7Z8gqvborKVK7ZI2jSCEHmb
96efSJqkk6rHU+wrIxffVVKx8AoxMLq9FdhlGn/F5by+BrzspWnbXIhFPqeSdi+MRLYrpZDv+1RA
AbzhlvItNifajY2L5lnDvUuKUGZyEN0hBUbmKp90EyRbtQ1lfwNAZG2qfTbkBr5l8mtF8OPir9cu
y3TxEiD/pku+jLOLcpCh+6L3cTgAevFiS6avDJXO9f0T1+/R76cmwaoqWyMvxA8XT8fScgVa1Ei+
uWE73oA68JwCeLdHos+wsE30n+F0RXllRvXcC/1TPgMJimfH/5dTRcQBeCl2IdNPfTJKaFRBYYC3
ppaL5ZPu2AzmK+DNSdIK0BOqOiJSW40NMrwI4wmSHc1U74mO3FnI06VSHmocOmVpR+8LP3EcLKKc
4Q9dSBAgrmi6oLv4zC5b3or9DW1n/1BE/OjOMqm8mt2FVdhUnGBN1OdjA+miH6jpINuCk4ygiuBu
X403YTuX+aEDN3CZ47lqU/7bbyAVGnDotQJ7D2uHK/QpzB/zO/3Cr+SySVcOQA6vJPv9bQHi3Ro2
NtwJTDAw96pB9IU9h7vWwwt1X+b5yKg2JCzgSXeDBUQ1Fgc1qlEZ2Z29hkw04bwhN/ovvw9G3ALK
1uImgD33L38vueA0Qjf2M+yBOsdL8QO144hHXUmo0mWw5+XtnZdpYjeFGVbKWYjnT9qTkgBgCbj9
dgOuJ0qaZkiK9r3iN42g/IqTMJ9llsjtwZtCzEQuWCv89qeo+xYTnhlT+nLaBan5YrPRbM4X0fGK
ZKDQMh6dgTaV3VADBxIc0ms9Xozvhn8c8rBjcOAad6iy9k20dnmBeeqStNNAqtdmEuygOLsNrtzQ
GJyBrdMyjHNah3wdbKFIYhQIeqQ5TmaCq2yJWUenftSsGigGtW94UgJlgXDkLSNYNfkSHqxp4Lzt
AxqUkfcKtFWSBztsC0N0NAMPrwRVTEdRB1Nw7cvoYbBEOuviM172XIOi8Jdw5nV5AQZKjEjhs1yX
jQAz1TE6A9GBenwlzqKimy7VH4hA+8Om/S9Lqg6ghhPF19llLZ6JINKFts4EckRMZoZNm3KQw2xF
PwTRjbJu2t9Hw1AI9eF2zUNdeCD12yuaU3HCA9UPhXrW90biK/daFouQe8rAiudE134V4/WGF1Bq
z8622xDy9O7gdoTpxEE9B/VK1Lhqy2JNL46ObuPJshtT/Nl0ghCWuYk9DHX9hk5L8W9mM9jBgcE8
tgHX5aLMj4taTfYr/Lh+7mgLklcCUCCK41yy7ylHmcD6Zktc23mfuMi8VuLqiu12PWf1j8zZS0om
rpgQYUfZeqSt/3wfetn5ySmTq+jts58UJkBCZuliF3eD+Vu0K3u+ifGetWqnBP23jsK6wdNbODTL
17qlaaU5K54YozGG8/nYuqf49aPHzyezzQpOzHtiVBnk5kBR/zI+922E/CMhX5WNHxzijCHl5tBJ
InUakAqpSe/9SSDl7SKsKpv3/IuqNWR5Jca6RWSjIYX6dZ6FWxr8dj3+/W2VPY9jSJcmRFdNVNEa
TDAbUi3yp5jo9zgHwWvk+0twFIrtrp4ZAf6a27XfLy8lo2Ak1al5SqzZ2x48T2Kx8RRUftfY+zXZ
/D26LB2jUKQ5CtkVwPe8f4AOBeMz8SdXptn/S6kM0+FR+RLyJqsgQEWV65jfW+/HF6HfaSbbaHNG
UjcuI8/Cydk86AdKViOzpZzFPW53Gs7ZdBQlvIswhZERzHS9kbr574Rjv8ZSK4GN57gUsg/3e2bt
yEY6gKcIsLR03AcFZMnBVj5XThXUJbJ3dpnvK7QnLCMoj9WfZwZopazCK8eA1uCsos8a4FxYvNZb
jO0Q5MmJf3+NcXc30ljeIomu2r1a+nbV2pnrbIdnV3hf8Hk7vrf504OIf1yGlepOr/u0qsQbkBmQ
xokAfrUlP3y1sl7Z9NGac6sQGqinhxPKxrUmJEFAUvtmdKf/s2FXMN36LsvIi0wodCCrrs0yq68A
QC2LVCvM8iV92S4Kvl0esOIL81A1GOKJxMAVqeaLC49gnVCMYe6f7zoG3HdON4PU47AhoyIiogNa
tOVDXUSucOCNWyUG6z+eFwQ3oy90tZHyR6rJL4tTJ6Yy/DmWFwvXsjRhKZ+GatoPPrFA3u1I3G/f
kqZQbKCWGVt4mN+clDR7RlKIffkn4/TZyLDZdOk0K2e1BeR39//OhqImBy7GzQY3p8Om4dptMYgb
wt+KhcfnupGA/Kh9IXdZCEB5nTtRSAhGnN77htLyS0b3ajA3vaUp6JY/Z6I4QrO2VLG8pD5KTJbH
Skh24z7PbLkrhk5wIimsGQ+C1H1ZYf8sQ6d7Nv3AwBOqovbVR7hvhDuz1GRAHjx8i1YfrWK5ImkQ
P68PjWK8bCSnkECM/EfxxpMuFQTCITLyhU0/tfnS8k1KGQL5R/BpDd7kEyrmobKJpLqqMJqtrZLy
NtvcxOzUtEQOGW/8YP5YYI2GZflFAmnlsqmktyGqjPxi8+z2DjZEzhrhp+EB+nb0IZjdFVSHP17r
7x09OHOcKGuRyyQIua8ILjh33nk0R+wA452ROYln74hnDC6l6C3nshaqoMSw2owYWC0xA1p8uLyv
mMVfSE+cyHd8twdWi5X4iMD+q+GVakEsN7tg1dRWMfPrnIPhcqk3ROGN/VWLi4gqXuDm68XKxaDl
XQse0d8JjoHEocJfhXhIfzpplWFteJYaNiGMGapJE2P4aqzxfWxgLLQoBMcWn3pCuCzgiUpcXqaP
hy6xHVfr02LlqkKCJqKkjuMjk8VN24XLxvvji4U9A3MQXjSsNgzadJ4VVBFf6QXaKVGgkUcsmYMP
42sNmacPFURSjRz6/k2LIPVJpwRbbmvmqd63ody0K5jjL8rh8vP/VdqVmEChUILJ9kfPAT8F4nAD
cjOHIN3DlU9ZBz+/k9X+50B8mYZCl4z5r66O0NXPYlU8jZjsZ10qFQMn5Rs7+7CVyst7ngWvFxMg
zGglDZA5sjnsfTPlo/nf0frvD6ehaC1t3VIOMcY0LzIRSXP+bmodtwdNfRoAL+/7nZpA0ls8g6HW
FY+n8PzRpTpAYm+0gv6ZTfSYGsrYCEIsu2Q6ZZV/F6db63QOLxDs7L6vN7Ajv5WpfedJdowPGNXc
A98S8uPdE0aBrya73CF55q4f7lBD8IeItiIPQ0A3nXWP/rLrrS1LZu1tlZwuQQ/yegWL8fMenlAw
LIcmO58T2Y6FTQU7OJiKp/MpvyQHi1uaKrHT1XFkG+FoVvwokPzebtTIlNip8BJ+WtmqaDw5irC0
Z8kXIc8Mo7pqTvDpUFzzscOpbD4MKBdDgTJlQZP1hzUItCQhBMdyn/cw5kxVvLGsPZlq3vbFYrR4
Us1KoD+W1L3WoYO9fzACv1mq8JwKNr8E8iX4EIgvz981m/tVcVqOHAQX/ZLvmwXmIHoifOPNweDn
ea1aExb+bjSv13+D47SHeHkpguDnzQ9K2HrSbg9rIUd6ET+h0GXYZGRSPX2ca6G9QUfJ8DIlKuY6
+eBjjYblb3ene5j/qhNfFceUZdv8UDISGugI+MEWiW2/hAo+Gtn+eBfnCnxuTz3ydnFg9j9BgYNj
Fsz+7IWTVK2960+7BXD+bIeBFXWcFGGHnSTuNGEa7Ha0/pFCzXKUSAEs5DdhbC4Z7fVdgubthgMp
8yQKuqtkXkUFAnP952ti5YNKxgLMDcFht+72ATl6vCi4cjJmICPPYZHGYVrpozDQwiDt8yjA3DGY
IdhRlI47Foc38h8OXW9IZ9xQFLExKgXiieQ8ioLCN1ehz2DgMny7GrhTODzARN/wQn1RlbrsNTOK
CosWr5QH/6Gv5XBGFNZrY78P6u1BOYbSwm9PFxPY7Omyy6x0z6y2++Rq/rTrddp6hulvzVT1RZW0
WUirDd/2ZjFpxTq1Ls/6zJiZxidGveXqfHAeDgGHexJxwL5CQa0wI5i9ausnI52pXXA8BAmlV20R
K5dxpqWU5OLfngvFPwkOrZiYAdCeSws9iG5zm87lFc9K06uZfn7rgGoknqpo+1QT21AidyTViU0p
tP0obldL5QCUeY9HvdWE9wXyGE5t/vnMg0Xl+5CroQY32fvHG5QjL+eEEN/Ue1Gp6/JmfcReSceG
/LzFn2WLzMqZV3r8kqIFzmpqnPdGwlwNTulGD7bZ32hGzcIvw0X3CraljcpgCPIFn1PSSgOouNHz
s5GClYvSjVZanjyZ7x++i8qtM58cxwcS4SxjQ1AGK7JTFrOatOvB1JFOJIqWoHJHYi1Unw2bMSVF
Z+bnnPdC24GqA0/A5UyX2ABaAQ7pUt0t/cUWABW6FtA5sCHdPVYtNqrapaixxoj93aXknYeDJl9r
OthIv1LkgH9spQxJI/AKi21W/1hVH9Wts8YLOOtr3uN6mtyy4/aLVpHp/pRYD8PBccN3hk5yOG/O
9PDPo3SLQ7JVzHLmxy//YYAAlutZ/ECrB1xdT1mp8L7BE3GyQZl6IY48+PwRX8h5j+eRFNLTaY1/
VawO1rvzUNVzGdxZ2z4mVV+YOYebXS7vNqoYMsDULFqbLkpclXNkwwjd7kq2zqa4bwSk7vNJfz+c
ysEuzEt6WqL2QHKW+YHgZX9wTa4IjCNyE/b2Ep0bUEvGgpPeHRcf9qaHGpPfaLAHpLzDfayMrNcE
LwPW0niR5sPZoUAcMlLKPvAGNaNyFboy9RH0YtHWlFbfiO7C2VnrVex58+R0MYj35ZIPu7bZdb9U
dzzZnymQ+AD2c8OQCYQMFGZtLDaegSCW1AXHb1SFKllEeEERjbv6wn2UWblyCuAXXVHNyfoIuvO3
f3a94vsslHCRwnOag5jw4BRLJF3WZvwB3l4aiwuK24UGvxLY+Q11Xvr5llNmhxc22wdqjAazYfFT
TbtbnaCHXnpmbk3C+mQvqo5UkrqtSo6zP1+Vt7dfHc6ZpKzzKtUnX/ojens/m0Wm1Oe2LFBOARE1
HDeBIKxNknDD9LzpISdexGyGShHbeU3IVpYOKUYJ/G108dCumm7DWYd08uSUG80ddjvlul9Sfnxj
y0UVvgqgcNgAFz+CxdPJXpTFebyTQnW5idQ7Q9V5lHa/WnOPRgrjYK+rgNpZTocO4FQyTGRNuNb/
v4asDa89EDFZQ0ySYF7yM/Pl38T+DfeDJD+xrTFrbrAxfxC58aPqaXEBR+l+e5jquKqjoBfYpZgq
zqnUavGlqiupzrZMp6SLFTZzHSPIXemimH9UfdTYip+zO53IeqmBsmaElKkl+gJuFyLBjnA2fGgr
GK6woGL0KfK9lxl4X93GuIcUPjJVB1Xlq1k3XwHs2eMxtYZTDjMNLNbYZmnqDBwHQwbp3B9D5g3J
UA6tjObZ6dpLwCtt+ChK8q5uukvohQvMzk1WfvUMk4QaVXVeaFKwaZXNPMw4lUKz0vBom1FFT0Vj
eQGrV8zjK5zh9jQXFwu6DswlMv+I/aaRqx5T2MFO4ELQ/KCpZOCI0EFaVMgmn/bMyHct5unxTWPB
Lf2OwRVuf19SmAt7aq8Jl0EmIDhD7UNBfCDDgP8ONwdyfmGQW4vGPgH/m8cu0YMBJI9EaqiqB8FO
0JUTjv1EdSzO/dz1E2tlSgDHJi0G4z5I6bAFnU9YEx0toKxXiKU2ARpWHxdkABbEB8AOVf90HMGz
8UMxSy/FizjQaT+4dRdq1lBIGqC/jDFig3lGN2GnW+vvKY6FqWLilwxKoRCZPSmzzcSCRxUfoirv
BOv9jRRD+4KKQCtje+HuBTCdyiA1+l7c9rsjziL/ugiQpQfUS9GqFEqB1d+yq2Ik1UjzXm5VEUgI
Ww/tXw/9mjUEh8yz5vq6k4w8820QIk+d/q7tqR+yaIjxqVvJZVDLIjwb2LA85uY2fH7bDx/617LR
Xyf7k/4ouvaQu1NsN5kGkJds47Q5Yue1lyVr6jXfwbkwIxO8iW48yo+laqoRWTb2RHKw+3q3mN7I
8JS7Gccwuc+zRaebr5VD0wZaaI5PrSTheBp9YTb4fswO4Dtq3k2HuJ6KSR8XDJovyGgDq1OsAh9U
WTLZjeFQ6d0uVZvajTuWjQq+1u/Do+l7K21pU15XjnVKezZyTA6vTTbzfeg0fiH6KB612I3IdGo9
AVmFoB+lT497tgXybDYReKtVE/nQ5VDv2SvKh11Hs/bhIoD0TdKn109PWAhzxh1WGuzX0yoC6M45
IRT8XDsu0gM54ogbgRfTHWFBB8ReaAogpGm+KyOWqUhRKdSNHJsh0a/YLosfip5clB9KutM+afiE
U3o1/yfra69uiW53w4YWzAOAVTGUawGMy0Pj9pUZPdSJFdX4aRqPQV0RiSma4cFFguZoIJwJrGfR
LpC7/WOl9jJK82sTF3DuPhioNU2YZ7W6dX++9OJvDLrYuFLlZiv8mqw3EHgjFaBRzAO89kydus7v
1lY/5ZZeHhVe/5EHno71rxlxR112h6PuxpZWBqKHEfYzimzSXcdW90PHvkK9dV1OuWHerQebnCCx
b5Gy7s8h6faygZ8ye2muuBmq5IX9ZeYI0ijBY2xsSkgxmKRQ67AHi8Nj4hIzfR+Fo+gLylCcLRzg
GxKQlhrXE7GT3R039jN8LNhhgaBgoKpgkjYRQGmWvx73qwVONPOpKbGaFrgZjnI+1xy5t6/xPhZQ
frU9RkpcduBXszZxzIUPt4pxTaG7zdXGedma0Z3em5802z3nBzgPfTe28zJ5zj+7Q5iQ9lHIeFLu
kvGfyMqcQtlYkOMESwSUaNpAjpijioI/hKKW96TUv4D8hRoH4px7BU5RvNMxRnRhvZGuH6z7ImPO
qJojR50Q7Zec0jax5GOxbHe6o+MIj62ksUvUWA+3IYR6oXlZ9FUP6Zb58YPLej1xC6ww7pO4dJJJ
jeRewbZwfMvTpSVT2TOUk3ajXzUVrB7cbyvA7TlNxRuBPhIhFQFGBM/AkdqTz6TkgZAgtEjRyAOA
3zea4HoO0zFA3ewLpOUNAHrJNUibBRtFUspfhkfVhSQdV9xQ5qAg/SUmya12kXdkGpTbZMpbaKXf
yboDzXRE2zXIPWcIwFBYw4xONW6lk7yucHkyCeNi52W3JtDe03z26Kf0WJGfR3qFsJ/9gtcty83Q
OqBmJXTxofJE2eFIvhUWsGbdHxK5N0IfX2mW1Qj2P4/MOYRWl9Ko9XFSc/9uRRqYFgQAsJqOKEOP
mPG52V0rTBYdhM1BKwR/a1beEuDcN22Z4iUvgaHE3JIAC9uCssS9ZM96wQhdQzKuvRWe5FP4HB74
1RgGQ4axfAl+4Gwdef3kPxbGs4iehFNDDu8iUjbN8e4ATr7AY0uvpE9BEpkIEePwt5Arz+XwRVav
5o+MWqT7AbYm5ycoybgwTD3LDACYOhnTXImmLracZJ5s6XUU668GhXiHrcqMFvvCQhzTQ6RnwIzw
cRamIznpY6XkpTj8MX0JUovmXjQCku2SwgMxRsU/eAnXwMdZA8tnUZP/anHcIriPP48iANvVESQQ
G4mZpok79xBU5IuAI7y0LHcnctGY8MylLnvi5riA+nalGoisri38b2VPUmOKTtH2c6BAXxZdpqt9
Ugm5SBsdjYLrdO0H6WHMhaQ/rilrKdCDtxGagSd7uvtzusFkAzi3P6Ebh3D34XJTsRcsSLCgxugW
6y/5DOPZYXbKBxohhWvqRviNxwjJNe8GdPeiYDE2ccTVWkKzeDEzeQ3yLhOCgc/9ki0kKX2N8i2c
jZv1M44ARSurqoWMD51bAs3yavHhJUxkHLCqyYJUc0fHOyMDj+Ka9ZJLlatEldMDAiXw17STI1VC
HBgm4m4DrXCopSOiMUnjNF7zuabiffE/1KFMJRcI2Pdd23EEBwtYHOX7q9rXISTySqhUbWqy0l3S
TfWm19wX/AEGxjywtMtuXXBQp24LL0nqLityojgQ9MyKpd+U7tekczn9w01/b7hGLAhptDBOd18W
X9aicsLqfBwsUahsJOmqLk5crj+cdSuiKTU3QZhQerYmMmyRJ0EZWCE4tWSADulS7v9TPjno1rKz
G/YaJPmtkIaGldHqohmfWgzj24eCmwzqmDj2Xfi8j6VLMYoKVd9x5AUCd2hZZ1lNYKcvIjqsbJAc
TauaFhYFmbFVGgKCA4u9HwEXRqwEJ0Gh9+5gBOyCaIYMTra3zJ3VqbJSc5e5D0KSk2ttQrytkmHw
TCY2d7Lr41tpJLObUVck/mxY0oYm4XSzvMRqr/chFrQacEeLSxwlN0AST48xxoUosE3k3AIjP6cY
V+pz0v/L6JZUebT2A4WDSxxqskkOx2PrkZn+1GI+1+tSsp96rr+xm9UayQvLz3gJr6l46tWQKwB3
jtdW253zmxUfmvuGB6yyuXAwz0Dkoh+xCOTNoA/Jwj4LcjfBpZfDtI0Aj8dLS/GsrHoOEWKnwAv9
ZF5ZFQuTq+9YMCgaAF/QkCAIZ0sQtCZjVzg39QcPBh7nMdS09S/G0wjHlOnKLFQcOysgMyAPdp9p
8maE3azSIAfRo1AYTKlESubWmVvlUrw57NKqiIEJyvtjcvFiLmiaNUsyImVs+oRJxWmC+sKZYcTD
lNVst3P2waE+75SxwlVOglX4mmhE+oWok3nVB1kU1M6tjh0d6v3deddDUpThrGEfOapEKe7kKUad
+emnOSFcbkDA4NTsGIo3NAodcIAvIdMhM9gQ2+MGLA6btyI8xb9JuEaICCQnBwGEmZPoTOn0O/Ff
tTNo5j0BRJCa+a0Gt3miY6XJXfUjIn80cNEDLEkSUlRbgGDNlX/uDwSmMCPaSA1zhS2oG0SqH8e1
J+JCxckFK+oTYe+yqBeJKNC6ikzeQJeUmMQFuNqgwYppWwPQM6lKgKWbiYw+3rlwzKYUTV+xrdWm
kxvnFq7cdFE4R8tsUCAAACiRYEEOSflqMVQ01GIFlzLdetzOFI7eds45nI7WXSb/kpUigeWfRjlE
FemZwP7OUXwb7+m632Kxpb2BZ/DuHdLhe6dta0upAg4iGaamGkQk16/TlQU6iS0nvId/IupPxDMk
6cLi18UyAhLwWfgF3UHoGXM5GgH6GF7qlWBhzkM8Gk/KN0FP6cqS4IEzWY0QVVZnGCsU67dYq6T7
hkrcxBaERVlvoNZF8EUz7nuUxGiDgLbo8sodjwSacvyA+VTOobAgep15toX6ku2VGyp4/am4KOWD
TAcPBdxnGl24rggXQW7SoC4aeGU0D4c6C03mu6/hYqgkDP5wZpptUa8C5X13HKpvMXZ+yxD4Efuo
E5LPHHGmuI7ApfxKRx3OIdGa9Bm6XjzwSIQbc44OEj878CalufqvSsYsgNfAibzLXEPxw44H4UO3
sRiYy4sXdJsOZy6V4rOfJQMHU2blHJPlOc5LQMrrPXmkZqsFEzR8ffBNhZaCuVzmuaD2nkyuK23w
ccJFkR/W/E6j8dLwU0ci+jOrDL1JKRY5ec35ksFABlEUlhYaeapbyQCK1lW7FftzSzgQFoTrQEBR
XVh0frc6hjiPbixA0SCCTOaY6srFQ3drzWkGLa9bHhfz69N2M1yTs9gRy/NtsgNxWWUk92t/0Gc3
6oB1p2/6lsRymyriYyU2XpacPd4CUrCrLPJP6Uhq7Z4Q/vFzW9QJbSvsUgklIgw4QAdwaLeypU/R
kPM0mK0n0wGSUxgcEI9iyHKbvJZjW8v1SwhI7NJDCk1gLC5RfUnbtPsNe/ByiKXljE9/F4H+JKJ/
22HgSs8nA0OqfVjPppkDbSUemhUnJudDOPAjv+zX69b5dhcjkghDqMqNkQ+EC9i08yR3KIz5ZXqD
nJr61JjIZbMQ0heU652WeJ94wMGfOy/ek5Lofmgtj0Fm3YqyZdXu158rAsZBiPUPPEz69BlOk0k8
bOFUxL/aGOsRQ8hy1aPF2LxoMqrfkUVcML2bmucvs3jOg5bzfq8mb6tu1ryaOBZz86oRD7WUoRZu
Lo0TLsOoXfI34Zc1P3OG+73anZNHXrtcPS2OCUmtAr44vxU/DYoBcl9FLVcQLr3ovrcByd9X9AvC
KNIRwKZKVS84cj0TNboGsSNH6xQbyjfKH33XI2z15lhdX6nmW+iDn4f+Vbi08l+DbdTzT8bsyA6H
3opxMRoyMCrwJM6oy3eqo2HAyDJR5BQzIYxt7f7tv5itnNqFyXurUXUv9LRg2fRd+pB/WLReOUrt
ObqjL7Rv9faHAlQS04y0OyP8CTg0MiigqfCcqWm4K+aL8UYf2OtLYr/QUBPitLZMtF+Vb2Xcvmrm
CG4IKU0fLLAS/yZZMA6tsUflYK6yMZQjIjpeaaPHX/vj6Ro3hGS0+85up01ym2NcRpEdwUcFKbnB
twzPnPw/M/lMyq/68NGeMK6hu34Ranyo/MBJlHeI0I/P7nHtiuGa/rtr5HTUDzOGwKsLQf36seqz
tP4tlcxqTt9fybkMBITnksnvLv3n7igpJPjncH89NIYbDW8aG+UD206ys6q9eQ1/YlW8NGW5yG6Y
87Lf11i5b1wacNySDZOYPFETvWkJoAZGbQhfnKyGppjaZPqlVOruTH2VJP1RGqtgBFUD6szC/9rv
ILZf2zZl32PG7zxvvEb85cogQMvsi7cZ62rMx8ndngqeV/pclm0ySyzH7VRC54lH9DAT+2VWgOl6
OrK4KpCJSbVlMcMXQoiUNrbF6Lx8KihBRzKc52cSUjjuG3rgGXF+SzwfLsJ4SGblUvAbQAuQS7aj
Z2luQErajogDVPd8kU019/o24zyRl+Mx/YOyTaDCwEO0vNGHFwT3ZSky4CJ4yFf9v/i3/u3y8/yG
TXgZOvvp3+A8UcNgTB88xaDJZaN9boWMTmcaEISCB9d4KVOzU272xDEsx2ONLpFtflUWxQcfxfok
liPFDO1FDD1yrfBMMxHOpZdNIMuw4F/ECt9Ca8ObxKisyrfKXBDDKoAmlUej5pHFbEwSZ/SoOPc8
rfBgnsyyG0zJNi76MslUifoTDJf8fCovIfxWLoqMJKzf2Jx13/AT9qbI3zlDTOKPOCCdT1qrXNJc
28ngdWnKgD3zoIe3z9lQ5tl0Maxx/odvZoHSGms5bz4Occ90XRXFrGyT9IxcEX6oYaYj9nRNUrPV
6E8VLLlp7a4S/As7vMKkD9BTI8qUSQ4LE2vzW5PFTrqN69tvOmfclolhi5hrvwirQPvZvsbPjcWq
X5X7bWkHAMx9dYWuPjd05m78nmoYNiA1eXXOxRKkzc39ydxQmX7y9lTATsRPhnd9asrSsS48enwm
hStxhhBPNo0aCvvvOV8XoXD7adrCebNqplo/BvETg6hEJC7JoWS7EIvsZRkaQ7uVDMlHl/wzuoW2
CjO6UfsOU6hX7+5AdjS36RJQKd2hImaOv4v2cNOTeXS3LuGe04H+ut+xh2Enx90RcqVfC3EYw/8m
Sx1rCnNbsYPO2fTPBj6vj5F3sePLlgOZlzB63f37LoNxVE5k012GUeaJBoV8bRwHrKOrK88Sb8jn
l48L4FU+svs2Ez4P1cLWkbPxbLX+tEUs447O/iZ8jX86luAozMO5neuV22xR/vm1GQOi7YES6HAn
jJoKtCg5ro6YwShqj1EDXXYtsba76n39/OhK4ihrlgRBMXsyRaAJ6wavFQREX7N+gXFX7RG3BTaF
FuqyOVgBjh9SMryixgx8FaK1TzLkPbhlGLJyh5HA4aSIJW5PzWzwVooTl/3ww2g264bScfJJyRGK
Ws7ZtwRKsZAee1JKSOiMGxWpMpTwU+U05o4N/ZXngeHRKgCbdh0mlJwNj1rKyAOhJpCFzcfeFi4J
iO83FSBd+zmtdHZs0ZdRr/NdVqOPjDZHVMSzFJhPiP3Y93yg9gqy4TI4xpKkHTm1YmPR0Yh8LScu
I1JICpUo6BYjNNtjZPbAhYBVbo6FsEByfsCgCg0ZXpZDt1i8vl8okz62nbzm2fV5sG7WMBm2z7Y4
kdpRkoBc5avhomv0gZH9Jv6eCnNS/eE8iiYXSwraxaYuuzqGGf4p2cMfc6YNhtfVz2wZTA3NGHPZ
PDxWSJYP14RDpX+t9D9mXx07/yFkOQ7dxp0ZN8bli1nUVU2YJbJvHd6KssyNqwPcVIIzyGnMqt4E
EsyfrKzDT4Wjnf2i5cM6X5BNTszOSRJL3BIpHptcPIr578ytZkj9mueinv8WSyunpGvVwy3lEYwj
dz7dk2ByMjIIKCE0lrfFl8QB+39jubrnW6+2Tav4VE6TEVM5YPRubMzuwGDUPz0C3GNepOOzV1jl
gWAvHH9Ymp9NQdsyD25o/CuzSdmpArY0/BVH+IYSkguLe2l2tuKhO4AYbA4w3iJq06SG271axEsH
Tldx9XuMAofgQFzA9TCCbLztOpxr9vcdbCq8kgiMSeX2batxFvQpQt+lpS2fpTaVQJuLrC37iw+D
PQxv7OE5np7X7u4y9aHMa5eSyn53kiTXzHGwl9Yp0CKP+rpmh8y1zqtKoqC+KcZq29QPfI+r9T2b
thzAHkoICXbRZECrelW73FKOBV06i40D38jpSB8sNk0XDjU77fhTvLzdjNr1d3/TJZkL84LodvIB
YyknmE/ppuKQuL1JPRhhAQsWa7NMdmjDg5W2cXzoEQ56Daq2zb0dHo+Vn6gwMs3GNeEu2pO9IvTJ
1lJ2sQ8T3s/EZBRDAWmw3bVIwLjenhqIkLHez0mfSfQomjjBrqON4i2aC8arC+rMZhjO398YcQF+
roSN3FKjULfU8vuw1QpOIZa1HJhNW5lOgrCffZAO5xAAWJpK1cT/rzyPttAnpey++EnRVuPTLpF5
edSKUvQ529pidw6Bb1crpAeO/oxMHP4V56GI4iUTWxYjJEfhAUXOIw7WYhgLkx5g18a3Vs0HJ06j
n3dBKQ43COcaSXPxUGIUTibW/uSo2sEvOQdRhdshSJsg/8K/DzglibxuHx643jaPV+c/TrM9eR2b
W/jz628osrke+3ZJmJS8jn9HX/P5ig7Aig+4iOurBre6tFMQthSzxZbfHo5vov0Gr3zSN66q4ME9
TcEyLJpydJYrwyExcWGYBa6NZOUWhtwKI/GKAvp4t/R9rghy/vEoHUhBr4GPfFQUzkgqvAC/x5Oo
pXKwASdpKsscvQKS3ZwMygwCgXD1ycp35jRYBtshcv8QLCo53jppyFAEKtdJtNroon9uqSkFeggl
bdbZ6ND86wKsLk4EFkwScJeTAT8VPKu4aPGD9s62n0EjIw3hShWKUnhTQ2X44/Zfkgq6Ez9TbDys
BTp8sqddhz7TFOyc9lPcTROkoKfgFBzQbx7K4Kb6MGiztJS1RaeITs1H+4C0/SsLJcFDJU/LIHUf
Fsk5Ou42vuB/ezBzw3Z2bxve8y/wn7RXJeq+5B+Ki2pR0UzhyG0sBNCf1dHWel/CJSKRSAywVYTi
C1+t5UkzZLYqfKQgfURAsUYgSeZ/IAUJBQ2prv7AyUi+aVqXDHzUbCCWIDZtxyb1drYO/wKww5kf
03ZgkuzlIAT0bb9XrvP5AGekiPKRgnBKUwhVq54jsOKguVDJisSMS1yKeCAVAgyMotRwOTDj7yN7
I1cI6qDR9iYeJpc58eaGguVbolD2SYbgNhyTqFMuPXDPxjEgJtnFVoMyVyw18yKj3uNY6RN+4/pA
vFiJWyIQqKCsh5a5vCDe+agWso3/26iZE+nxves8vxVJb2GOUNPssK76wvfPd9SV9JEUu7j2f/32
ca1xrp8tEV7D07fqgDqPcX/RnJXxNFtzFSHw8ypB7PaQJg7a7r+se3ZPNOJQ7+KQ9uhnyFNH6Yd3
hnY6r4ULcGHnVZvgZwg9RH5Byixq+krmIvPDxpXJprdmj0LO32oV9cfkGhnMZ0abRknFmrlxHFWh
KXH6IVVLIfVmqh++auYmoPU+duZt9EKHjTfWL5QtwwuchNuwSunWKGE9WaGHz9mREeg6h1t+tiyV
UZc1RbynHNAdcAKS2puqh+4gBZTxhaIyxNaNyExx6DaJTOY20NAFJwRqWYgo/Nte+4WPD3CSrcL/
gjm5rmuXGjWXW8wp8LrlZ3wUnBiy/sREaEBVO8o9yQJrPFypPrEfj5US0nmw4Yr7iq6FaMk2D1Bf
Kdn/dwsgFjs9/X/u7dgDl+3re6efOose1GcyIHF1MsHxt493Ee1jmtjN6JhZCPDst8Um56h/PpV8
P4EQ3dijQ4vSZhn61tyTX3pQ5gWLTDYYKHaMJwE3VAwN3YtfN5eo0y43p9nU8r+DbvgUMuPqEsEZ
j40I4R4wWxhaIUNtgy9OHjdg7KOYNkX7fBZx7A7+wRhmvWl4pxVEmChROdSVmkahdw4kPebcDH7D
QkNxoaMc3nfi+bB8C1oq/YSsYnhOlBjWu6NPv44nLRqVz5FQzscdyKmHNhGOjOx6Opu/V3yVBAKS
tIQ14kHUxD1a8Gso2eJW+flXUOQ+zjuX+evZd8t5IbLmXuCAuRBzs7urWmLcfthaoOCPGn/6CdAG
E43zDjg2q5oYmoVZdgwwojEskiqeygpH+gLaZXhJtUH84tvtn4neVQmBW8fmh3Wi94wSPCmsoevi
zgZtO6HykP9l6OqKkN7zeGFGFo9Q+tPcOa3WbAEP2PTEDCXpLhyUIurMFeZtdBuFGOefgPjyhHvX
3KUjuCuW41HnrhFO+786nKzdxcZDymtw44aBo4mMUIgzzhsKUP327BvgbyTejQXow+ve4f1HsRSO
F8tlqVddRponk9LlRS3zqNUPYcUPQaN9f3h2g72PidGFPcsNiUTGomHXyswMdrQmC+hYkdLU0Iub
PXUfUMy7Yn0be+b3w7i1jmO6UmgZAWAb+fZRgao24Xd2DNzWhpSrDbJRPdIHKsHTdc0BwDLoRIE9
F6R6DPJ64J+75YadV2Buf5Fwog6ux1+DRBM2hAi2qed9d3xjrA/9pivz/tWk6UV84+sO1TakVTQk
PrT58jKcxdEQptE31EfrVyIEap9guxV7Fl+/pynO3NzDb3Ya8cNvY6Nn+VB2bqRxDkAAJcshy5zM
42vxikcodi67mGYcB9ziv7f19H6jgk8uJ2+quyG1343n7qrBFkE8CIDRtNtfovVRaPPJnhsKJXmP
AuPwIZPb8y7Ket1MSktCJn8bTWcT8vBiXM+tNHQ3pYV3rBOk9F7FJi1km9ye1s/zhYDOB9xbkcYw
ENmAPsueNAU+efn1xE5LCQGBxzDHD/K+obWvOxLhuwYr8nXvLhQ6M4ePA4T9X8aEGB2gst/Wnzk4
c1n3CtyPZB35sFMgDLa2sbPd/h70koFFN3rjMyT7Yf77g/jbDTPtdecxKqp1Lr6qnK+3ZF4aDN1d
O21Offo7JyGOuPANedPRww7e2P/7kA8s8YxuWcmJ1TqFo38ksgkODl0vo1IMYvW4UxAm5TwC2PEz
Yv38FV5oKwQ22kFx9DtDkFWVV3Wxj91TOUaIpsmXhfk3cY1pKyswJ1YE7Q8q4g9+uG/BTKZaURvo
IhHX0p3DBSaqAQ0atNHg9SZiuWFcCs8TI6vA+EikKo8yv6VrGUm1BhlnJeyLSCvr5QFABvOTq4R5
SgaYOYTisMSW1F+gikQojK5x51+vlH5XT/iq6X1oNmzXf+jf5PqEgHkXPcYD0R4sh6/tsWWsCkks
wwbff+aB1ODub6qFQu96zLQwIa3vUTwWsT7cv7ga1IZybtjYZXsk+vuzowK2O4OzkPO+ILwBYy6i
/3/cTIVhRD6k9uuHovSW1kWZe/yECqhl0rxd1ZqEb/mIOR/Vn2TdpWInv3THyHoRWraPM2LLxPTD
7Jg9CHYj/koyw6KmIemO0m0vfdwiH7733Q6EdgXTIHDJb1I0l2S8POCXepmyAYHC8bj6aQUw/iA7
dbOQ/Xoa78iZfmfSV9LEC7U0wm8seQ+V/n890niqTBX2yVC7qLDZR/qrc8OcSkpAzpnNtFmOFNBT
lE5l4ESpINkL4/WD9+0FEzo01LJJ6qzmoU2AutxRwDsd/DsjIj/7eIYE3YIEaUTtPJOsnxVWvcog
qSqkAWOKQ7gsoQ4aKTzEuQMjiC4AFK2ma5NSlT2kfS2NftTQmyoh7y+hp/lIgxGKnLDWkn5Tk6M/
Jejn9GTnX7kQm4It2/B7FmT3eetA39dz6Q6nL4BL0eUhqHzbRj0KEWmhgjPcUUbsH7c/qrhJk02x
Fn9Tb2ydLNNNySiK5MmQkNVpQpk53gSL/ut1kCpDU6Utq5BBjuKievfoAhRGG43jXWVNNK6nPs8A
Z8zBwqFmmuJ4ZuZ92HFcPQscdpTXc0BWgZ/s1Wm+nKFZyS2uES+HwxNgYdrrTrnhiOBGcwifE5V7
SgH/LH+tAS4NkKmf6ap00AzW9/Jn/pGAD1mODGzcGpYcrRuw3L/oHj6uYJQX4dKDg4xbU8DDLac0
fyGO69klUw73Q/Iu1ZAiLtYJ38l1lIoMOg9A8Aa9QTgOB1w8JdeZCyaxLiwrGT8QlzPIpwDT2SoC
+zloCd+BgsHzTVrYH7DGoaix6BM9OeY5ix8R1wyj6Ag4mOY4jmftyChmPqC3jHBMwQD0ZbdyBq6w
GtEW48vE43qz0/o6ftKS4xCVw7ePsyJX9CkgljGCbfNPdLicloLaW15HNiqXCGzhaLVaalyRyKpR
gGKANrx56vOufmwOisivGqVO2DxI+jfNdTUb7WJx1A5cdhUVQV+E4a8eKhcbqhwypQdqPCYIfmnb
KsHi3ymI2MFF23sipZSROLMbIR+0hZFg+g0L0IMkGXyn54+SaRHBQgG1Xspw7Gm4ggwzSaPpG8nM
fOg0JsAKX/6NJEiGUpCC/dPtt6wrPtAjV6N1Nt6XHC2txD+CezvCe6UB3K2VHC0v4g6LMDV8nQJl
bOShtxjyLGfmgp8CP/mbEcT06S5/2N9KNklzyAyzoxoFBy5szjoPAeZ5dGYxZu5qRk5mhKj0GFfv
RUMgwnnQC5EgDbOQ6RZCp5WiQC0XywUVr59ZeFsnV4f4YkjSrZ5qlrBxyXIN1KTJx/QgPGEeizlK
z73JIdFDO1wOMgtMunhLwTLWOqVeDXrb9Gu5wMK9g/gAKb3+V0yWi0efkURJjVnU+TPRFmg3SntA
AHGPFqE3FYB1JptbFojhCBtumKdrUgGpqEjVpfQRU62I7WCL7PKgZJ6Rz4Hv6cZSc5r3lWDe7zKe
VhQV6X9gYQr0lKhEFDQ0ZVIW5yfDE+0VDFTB4Gn5IxdO8wRscyookAphOV4Mexhc8Oz8pBubYfoH
0IjwxZ3MjryPva56V43lLNBDR363Fv1pczFa6TUXIto4t8s4FBsjiIasjWYKFQMBb5uT7ZQZDiXs
a2WGtAz8UuC0D7p3yXjOwLytMbmGfKqd8QXxPtzcdz7YIJ3ur7B0MsWZ8gtfkiOCdrL531gM+w8O
Bb6gRhwMTsVC0TyQpKYl6wK2NSOZDOugAPFtOEDGj96KK7+O+tM2oqy+A7Rx4G/XgtQ3O778IPAi
tbLA8591dDJj0LASOLCP71Wk2aVC9S2qz89O+FWhUmDE1gzvS/A3NmnuUqGLDWXQdbQyAO8axz82
zu8PUOHsEtYyz9iOM7g3QScLcZ/mEXGiEwLjijPj3TV8hLKWp1u4P8UB2iwVoGSU2oynJOsn/ezT
1VLR6G3v0tI0NqLCDVnz42yvKURtKnxoLK0unBfgp/d/AuAnrHmB9NhhR+enOUswkmprwSGxmqf2
FQ2f3vfi5vejzKyxhsEJ4nnWUHcilcQyZSnjVLua8rT7JNuRIkp5LlP1uA6APfURH+ue8hoUxbLD
a9K9rH79WOMwz5HwQvyy8Ix3jonW1Zm2E4fBPTPRMhmKRR9c2tp3dfV3RdweE5xNoZsQSamCCKz8
h65L0wkFr+IQh2MLNWMu50A/B1Ohn65NsAUse+tOiQ3rDS5oaTLZwvSZts4dj5/IemcLb7NQsBC4
M14MZLE0q4DFrvFAyRRIhKe+3q4XLfvNaJJqspCP0mBr0EkKxNN9QtyeEV6IwnJoOF5rgQ0maWii
0VLhX9ILY1xZmvo10Wjk6bCs31YYRTVKpr0DBUMXGp8wlGOTkosuLejGQsbEEVZ1IPGdcmEeNJmT
O/zz9/9h1dxKhsmh+0HIxG6r6i0sAYnbu96owJSXLsfWiuktmfxtI4zjvgVIyseXrQSXOWAZoW5X
oNW2ea/cRb/llBQaj+hOl6T15hHPkE9xh+llgRtYhb/HSlurDGX7jhFJuWrZoc5vTk/nZrzW9Fk0
2za7XzhgMgtpgf022g4J1v2ZUEjGsmeLNL5QSX3Q1etDu9td5y35xlorszIt0m8vdK0h6sEAu11I
d8I+3IEdGKxqPv6u1E8NEAZ2NodXF0a3okK7zgiqHda8am3FnUhqjy4RXYhNmShjD2EWMP5dEhNA
R9gOrpudMGo70s7Py7qkah+3uXazQekK67wdcnsMiikuFZ7eOeb9MGskQhZDoPFYX0BJmYwrUPWf
smzFM6px2B6qPFaCdO3Fn22J1lx7s+FcYpVaDeKUifZpnk1VM0VPrf4fsTNct8dHNVX/ntwhwpuJ
v/6OAcSSQnOH3Hw3E7bxj16tF8oH6boj2U/xDZ+pH6UQOaofOjd/vHvviIJ4sxUHy8beXGMLMlh0
fHRg8ntJ7ZLuLKM1QgA2IMwZ6DBOqIm87XLzWOyek42+kk8x3/G99EAkUcJVKadVlL5utqGy67Nx
O+QXa5bgRgnkGkOiPOtKw+spvSG7ZOtcxeSkY2U4GfJEyCO27L7095+WFP3kNdB/yT1laWRQiyFY
EL739C4cOptcW+KYbO/843aTbk3U2hfRDKZ+xb3gSZth0U/bjtBzmWwHbkI3DpkCqYCN8yglrs6Q
CMDLhB4W4ErrmOYEYG3PxKOxyNgFYgJkpjhwth3QKMhXYbnRX7J3xUghnP5qIzDCJICVgrTgaEgy
r1GPmz3upt38p7rmozfPdRAy/pGrk+Jsd9UClAPr9Fw59ymeVnLCiIfiwDN/HVw2FBXc5iWmTw68
/giklDOWv7vAI1LRt+enPNN18g2NW3hSqwsZgPVGdUryzxEqGMUiXoydIYvt04JoBghTs6yHckun
crr6tW0PQOhB+2L/CUJSmp48/Xu7l6zGp5c40kAGqUyYroBqqPXpHXDibsaGIuLDaMmGDOZMjqb2
k65KwzC+X26UsuimieWRaSaPKqfoKP1r5YnhrCeHJh6JXmYWJSPWawZ6FNIRdzTNu9Fljzd2rorr
1zoMl4sHImR7SbP71C6UgneF5qfa0Mh6GcKJNwS+Yy0tfj7KKaVnx7rPuMLOt7a1WKP0sMoVifZN
+bucYLM/fVRlm5JHrW4PHwc8A4Deh65G1/ZzA2wFPdyPowInuZPDpgL9ujZXIhFVGScP9tiUj9Z8
k2ysXWBMtp6tPjZh9AXOSnN+Ap52oTiXJ9TaRzGicd/VyHOIfkl/Uv6EhKtSZG+oqT9PsozUF1c1
3rHAXwCfaviLoGotLEPf/+W8bYPYP8XQWYvtZiriNNAK3lvp5MOu+QOruVgqJSTD3MvgLMGGLSnl
m3zWuIqYZfavRkTIcisG5Hasv0OqdSdCoKi4a5+Cx5KODxWLykcwayZ7cDOzqv31GctAIgKzFITM
pQ/sRCocDunQv1//8bErYJ6xTSE045X6Bw1CqNWdLUQ7BwD+gDsBDs+21LFHu3NQDdqofSKSFNxi
WsRY0N8BNLodFi55jx+zi7SKahQVxjkfmFhSbfGHEMCqjU0ej3HblzQocdI9DAiRUI/8KJcAMX8/
E7WuAWqXR1VIjkYXgrs7fi9COgHxOmxgYfTzHMXck8BkQcDbg6znZKA+MUrD+gtNxflm165bPCMU
DQpJHFwW57dvKNRqnZQmetsGIiQ3i24ZP3QjxQ0ZvP5YC8nE3fFJhB51jIP20g8brdAtYFrqW+9t
2W5CSsdbcj9wLIYLYXySwvaMRGnISlo0IrVnS0oEQ60HdRT3iL0KFVtR2/zE2vO2Zl/Ryx6hni/H
4ccRqDHiCae4qFMVdSkYtjBaQw9IbmQE6UOcNd5Mvm371aeJLMV6CmZSsIp2Ga2q+AhkEV0fvis8
SJDoO2/Kzl6+sHF6vx4hoPODYXFqp+g7wYNq6S5JZ3VB+yF3c9cLtZlW5hYntNNs5ktlD6gR0Ro+
hFjZdtJMvai59Eu3w4P54J2eBXpBvdXNvNVu5Zf5hUie45JsLGVhqVQuRljDTiJA9uiwa0XVkfhC
zBFm4ObSCzrrzsoR5s/Wkhhl6Fw9xbWkTensgteI1Lv/4q+usCcXzKr4ZzdHLXuV/hRs8oIeZUJJ
W4FQFDOLQNHhqddJ4hkQYIJ8TF7ft/ifcCQBuQFS50bjzf0trJaJArR+mOiY/+RiDGOcCSh6J3/M
3JvPtngqiDAN8hf7OcBdz8KRkK3Sod/ESz0lhrN8xcw5C0WLG8SMKsmCRC9qr8QlLLosn5k131rr
wc3ebTTrOYR7HS/weW/gmUa21M+5Utay3h9Sg1tVX6iO/jfmCj1INa+zwlQ+MHc7Gw8faWxvCgLc
nbKU3r/PyfMHJ+bvVzToZMtq4G/Iu/GnT+Okn5sy1yc1vkN1t+6cWcH7kxEuO9BcEL9fzDkeNbhD
5e48kOTBRy1LxDjcwlc44lvJDNLn4GjF4pe9HiFeAauIfGd9G19h5hMsaPxWTFez/VxnrLKbR9yk
hWyksDoFpQhZT6Ic+VAn+zGfyBwO8BoZETtwRjFwRdhkYrx876Cw0sov/TCVPWnFHRMhGNSZrM0T
hOS7nHd4FMZ/uINsuLAuTfR01GAnoQ4bVg6NJs0veoP7nKcXrK+6F4vUDf3tf+WhHuChcGbRUooH
5+z5FiamyImukqbTkRjbmMMPvcTe/sA1OX2cRVE70blP6b99+5btBdV7r5mVEU9NuRgTYbwEvz1B
UdW3TiGsouPvNuG3Y2T5mAOefXXLEuzADIW06S0PPJp5aR9bc4ZVUJxfwXHZ3PybvG+v71lUB5pq
hcu8aWDU803ODTKMGFng9ui7AXnf4peJ+kelUA5oyXw78O2Yh+R9eROYfiBJXOoKF/fXpCmANH27
dRBB1irFKapE9DatyAegFpvswtXXfs1g3HZEy1W6sAIUaOrlN6ZkjZ1CxdUKlEIlbwyYG8GjEqv+
mzwDCtFPUEP/39lxditOqU1LQR7Ev63xUgCuXHkIxaGW+IYEWem5geUbP6sWh8aR2Ny2mNLCkjbb
5y7F1LQ7wqgVLQ1zKWEEMq/MwAEJKSpY/Is2CcN6l+e9/CYw8trhdhiK0gK7FZfYUwJ/+zu/4QFr
hQkS/Y7EAP3xvfxi6V3jBAE8ug6SzbaYkkUlac8hTvU5RTxOy6MzyU60v9uDs3T8Xamj0ndTQvJ/
WnvD6nIQJxoKqIl1LFXJMH4Og0JlYJzpqcnnfpTN9MHdRe+l2wJlBtUaC+9yfkSxmuY3ZWylaruH
R5PHkycNQ7UKa7Q6qstF/mdSs9dWRbpV/O4k65Fm5QO7IxON19m4lCPKbmuWi1Aqx4WU9oFHVSIG
R9nZ8ul5AZzfMBXbWStQK8qUIzEkU4DWnU93MvdAPVNbpm6Ftn2qJxUh/10iURlZuaKgYVBQYEwj
9cETipOIcDqRjqYZGqldIIB9wTkYhooeY+Y01bso8Td0Cmim1/avt99Fj8+BK3ESpaQXBbW5VhF6
3HRDNQiTUxyYK9bHRU0tO5SnuJAcsvh21qQZvPYfp09xV98/xGUDZNBykuWrKd3DA4x3bmhqugGu
haJ3XgqO+A7WOHSfyVUsBwqquCJu9YB82Mxhvsi03Sz/v0neC6Apw1aE8VYzkSzSJIXEV/BpsFEv
PRiFq12FYjV+Yt9Cl3YSrlIA+bNw65wqv9+q9xTGwxuiM3DbG26ijg9RwWsfGNVgHLkXq5Yy2+So
9K7y4PSPQluyvY5GZW+e19fSFD2k1OKXx8ufn9R0LIP2LN1La3aCRo/mIAeA9ShFmie5s0kSOasq
Q5DiOvpA6oZK1NVclvZgnqBck9rzsDMwwyoqZ+Wn+EdvKYtxeHN2XUHQtFeRR2CdU+Dbedusl8Qi
K6hGr+MfZUZ5kNMbmLyDEnm4vnq0iaFZB/GiUacZrY1H1qqu5wvknRp4ciShaIdSrnGGKWEIsdO5
jNg9vufT3MmrmpZTX9aNpp3nsQS9XpU4k0w9a1tokQEmc8R9P9ZiyoCpCh4ov0i9GhcYEpN8TQGH
Yqc+M1KD0tn0rv+ZJlav1cl9jCwZkYNIvfFop4plBuZAvX27rtQzx9ycVU25hlphQBNfXJ5fp3Yt
pTc1gJVlzOgUW1AHczDCJOeevj1hu7w7qdhSIOcu3FuKjeFX03wFbcVRqZ/fpwbZuao+VH1vYXX6
OHqMKXU4Q1qA2eyX1RE+EPW3+L9EMu6Ubeba/9bI7VHvs6BU/vB4+e4M6eSXSYK9YZ9IVh6q4J7j
Vj9obrpuMBCtCzjnGutr8tjn/JyJf5FrIejJGvej0crIbq+Cm++Tvk1j6YOY0mOE5cu3AyScBRUH
KLdPLN6d2Q0ozjqtdACjaKyXW+VUMjmuO3dwLAmIEAIMv9kRfhtoq7j5MDeDSANAiAy5gYWVAEP9
8eeJGtbEHr1AWbcmPxo0E7TNZ6EjgR+qjwq+QXCxVnfGSDW+IR9tXZ4tU5Wr55/ZTdZlk7l3Y725
QII/szKBbjqOPn+A4goilDB5h1hjhFiv2sk92pK5cQvgR/arXKbdbqeSNrKElkM3azrdMV2bpYIw
rgdNjBHqI2VYpi5v3zyrAZ+niLnX4qWbfrqjgDCliMVAOVK4uOFhs3FICZ2QRjHQ6bsZR+RLAKdz
n412L4y7tWlGD48sSH5/sYbdyM+Grov/QkGXeDuDLPH+LzIRzM6OrzodUTzZN21T8PztrP6yS0Eo
N2jGLM908+UIgTMsqnpYYL/JMVr0JDeGzbcDuhW+xI39oQBiVYoNHpYAQXpDWHOv2U/N87jZ71A+
EPWSpz/JIeol2uCXj3IjtdEbvFblUD5g8Jd4nVhRE+vASS21g5pkJIWY3hF2u/WddiRoJ0NYupLk
h2GPsF60NL3daAWooaj230wtxGB1PBMnX0Vce1EfVca39Kjkh2/rtTDKN0dotEt0jCIZI+ygCNwB
AyD3J9ysQvCBVdBpyiUTzrR1ANPovelQa3qn9Pbty1Y+mBlEPPPTTp6hnEk10DH50JtM2+4ryYRG
3FjZknm0d1nLNU3a48KIBQUYSEyog5MiQSdWVv8TkHwAyjGWzmo4jHGzinjh3zL3BkvNPmea2fdS
NiymrxvDdduYZZjroxs1nzaFD2HCFposJz7FDVsH67BDGYOpU/aB71Lp5nFKxDHv/kJMThxKyj0E
zZsVPOs0hMAMhuLODJefHNfiqjBZsGlXab0xBOh1rhQrByadcTh/vThTcjzkyNCIQKJwPo6iBPQm
OGpD8zRYb7VsIQY1AXj4mLd+ZKSSned29y2uMpV5BVqkCDgi+1BJZZ1HxNAM65UAt6Q9TDDr/efe
9fq+/POoHJb8EuAqsuWPzA2Lse8vet4woun/ZopBuLhqWjatqR2rUXZaZYVcqX0kWMTidI1CWr1x
j1D3Opv/XXg/L5LtPh7Fr/QaYuzIVrqj9pIz+j3037+lIC8j8dwSlGtaM6+HB6q6Ar7tMZ5Nj4iM
nYIW4ALQ3fXMKIAL660qt2s3IsYNv+YxmTtkYK/m50VqVKPfqX/Su6FUNFRgGWiyTngyF2i+AiQh
0QHmpPGEPFjtB8rsXHg/lURVhJ7eT0d4QHr3rmRAWccGaHrneo0RhkJjnYulDVKQeVMD1jaeZHYi
iyeqQG2NuF2BHhPFv7bMCCQn9DTAv670pdeOsnV4rAML3rzGFLgYLIGi2iqxeg58UBt4PHMPeFi6
dDRejL7owg83S1YPdu1af81vUMgd1jkLy4bEMU7mYViHED9j6GxPOt3uR5fOG0YJaQbGyf1BNEkT
2xZneTxLCcobf57S/iJE28Va7XZcrRwxi83MxOrxR5kQdDk7nGThehdRnAwpw67QcFpgubcCFnQh
+wNNoDkikTwNnL9OBbNc8v0ou9wOKBLxVPa2j7cU/1MZlvwuGuHT5L1SMLb13S1WCbP4+XhZV0ww
4mB1WBf4ZwnFxe6HJc++R/tS6fTp/UrqimqgQJroXjM1aawXRzGRbDxQDkY2r88/VZrHb3jIBQKL
qwze72i+rDNIo1j9GxqgDX//er9KKyjivb4sA+oWPQjT3PduiIgQ3rMhdF17mZUwzMZsFS0eQrPc
o274dl2LXM8bWrcvdWpQ4jGpxLFENpUQui+nmDXM5Obn+eyf3iuaGsfLT5eE6AlsxKslZ3XrqIly
ZuS6WNQBs4iplnQvinn/9Au6A+W1tL7Wr4avKuWNUcVHZ+p9RmHsqRQL/JTQxap8ExFWgfHzA0wG
Y4XSCVoa00ctOAFtVjoU/cSg4xlM8GSYpNdJeNt8+BFASmas4bNo+v0TaErsTSJtIBoeiwwzcm+q
A8Nce7J0JqmmAt8btaAZ5OoJjw7hq2dOxIIHJTzKWvZe+zA3P3J84KdmruvHrd6dzi8aLax1GvRT
ZVM0FAPs0YA6cwL7+Lx7eKYI8eJ/QvR51z/yDz8CVQnJGm1Pyg3KSuKi4E47FSQyMzvMof7Fgf4B
EntphhVmPRa+hLvS9zCwI+CcAwpSKCkuVQjNn2o3E4UhOrxwARNXPd7K2TgjmdX16i38Q2dTKipO
iuFNgqKn6zUvhp5tAlt9cNqS00KXJ3IuyXWFZ+kyFIC2tyRn6vTEzvobLRNdWc45iRJwESBegBxe
r2ERWua07+aBaPPX5rJGjAoSk3NWom61mXvXLKXfVQQuldc7JMO+fBJguhNYQK8bggQgDeIrbquE
7eALj0Go7Tak74RzXLtfXojsxncdA9SxFA2IinM2dVhecyVsnCCqbHQDOFTDKq3ry+9inS4/K24X
3qoy0eIJCn/Q18P5BeDhzEOwEHPe0wHMc/Kd/OZC+JZvNjQJN6/1ipdHoUM1G6t2k4qSaYaJG93C
T7jFGfJsAjBxYb+USFVySpObx2+iQmPJhwUGY5tYKa/SHNCKsmn3kGpZCIuGOt2zgKSt8tYVP0iZ
SH7R7naM8QhxWSvyPPYL/Trkq0u8X0TxEXJV2UwHzNwctPQCbQPvktT9vsvcno5ntFIP7LJjlAiv
ZASGXupI3e0FHDOlqrf0ilFhXlJcEqFUXn9bDrd2m7BotjxJkneUEyeNBBA48JxiypLGf0NFd8C0
BUfx9cfpTYapcfjauOuw3HXsoZASe40JAKnEmf8XAgW4upD0ZxOG2xmntfcnDZr85+Qkmb/EVA6g
2AtDbh3jhj3kMdzpMYFUn84r69Q9gmOa2vsSRi/TB8KxYz32JHDDgcd+2dvA/GgnxOm00AcT+LuS
X4z5n+7/GlRSy3XYo7A5XVXKmHQR5PhFebGO1myTWpdj5iPK9NKNIseRaVMMNaWyMRUlt6FN36Eq
S8TsUT0sI8R6+wJ7RRAN41TkB5i0mUUUZEpqYgF5c3ma2uvzCrM9GVAZVZRsj8P4gDbA5ZOaSvLY
R+S09AlkcIBkCtg/ci+S+Ijhfm7AzM7y9PGR7+xfZDKDxqn6VaksJeG32z7wSoXIZJQ3qHcB10O3
QKu6wkx6mnm2FIQi0Y3uEfu5XBMSw2lm/RFgrA23ZPNgWA5CVyx6FvqstUb1adV4EzsHCKbewwys
vU6AcwHq1+qXoKah05LsELUsMkvz0kkgpkyFJTarHd5gkcts3wa1My0Pv1NPof1Ah9+530h8PjvQ
HKIOJwaRJyKygl4NDEs9k39ed8BCbRwiqQr4iiG0BSlNoB/4lyzvU3Ao64+jYMxyakhpo5x8xO6/
ufp8KEyan88If+hgEbxtrHm/CNaBGFwZFSPa3GvBEamKkoWSV5K2pPUY2waM/VSioSoNQtCs5j4G
XqQz1EgJfvFJ01Sa53aEsQ9clDTbxnx3Q937Gg6vy2aicdyrc0Qm/HVg9f816n25PRF9XL3Thft6
o8OcA1Cv/p8T9MHPXDgQWFNp0WUIVLwq8OXBwp6AVnYlgxEqi4WUGDgxNABijUVbireA6KiPzs1/
qSsHRjPVrSEYh+xBwzeZgL9eBkNu9gdlsCJzrnnLsLp3ydSQd5/j74fMvYE6rWVEaMsG4b+m7Qau
R3k4i4XQf3wnQT6n0XZ5s6ba9GKNhT3Yhn02F8S/5YyRPZ7xKVicOxyLai1w9+ISjd+8V/djRt92
Tt48BUPt9u0gXBuctYggxaV/V9gmf1WUOW1f4P6GaoyHE3c+34HwVnvxg875mq+tNfFcjCqZpUVU
L7I0BM2BjVLZMU0LozFcltegVby/4H2zHDvdDt8Lczu7b130vMyolGnsLPSmYpI4skfjwotzpBe6
2Ht7nqSpZRBTkGeM73MEMgO/12j5WiUuHTTKfuA/Uz6z/oF0z8pYI1XzuNzFu0IjOOGGHDBVIBpn
docDyXNWTl4rUJ15pgopcfA9rh5GbvLW18whc/uw9eoiymlO0vvAO6S6hIwcYrMdiz+2JidNdeTu
d9xmIXkKMrSKE4zko6Q+YwQTwifq4QVSN2oxLsbKoBoZTu5V6qYZTuhPCm+wRn5WYEkv2us7cSBI
B/mVnBsZ1NU9kuMxjoqgh5gdfJFtxiXs1XuaaWg8v3uFIzTa7+OEHCU9krmoZiQCcAzMS30zY+Jv
VewRDt6Arv0+2N0+JdhiEWtJc9kp+DCexv91/9bl4G9TRg4Xdid0tl+nCTAsxEXj+RotPb8UjZiM
MJAsEk9WLozUH9fKBFklQ5uMMW20x8LV6h5RNVsrESsI4BsZ6F8rWtUG2cjSm80ndU+4L17slJr5
+M64cV/C/s9O87bFJ1+aGjjpecI7GSfbkeIffS0Hi18iF5lTB/+hrLRRhMsojJXZZrb82a3RmQse
liZjclnEFF+7w/AyVa9IcdVsV0hkrvkdWzFI0Bjuy7yeF8JxmVpMRwu9jH3+kmYnk1Kjj+QCzLkL
w7Pbde1Qs7k3WUlt7P6urqx+piYqco4Y5At3BNUpXldK4i7HFZZkTj5gq0Zy9TZWIXm+x5CUcWQ/
LFysfkcQFtwZcT091qMuS8NrCT01JtxTHwPuPGLVZ139VeCM/odTmkK9Xhqfdq/wh9m5R35EK7FS
U/FplTga6rdoVc15geb/5dm9glwY2jp5h89AR5Pz4iZKpwizUTdja7Zj0NYAAW0q1hQRzUSBGCBf
LnYh5Ts5XSNnpqwh1Da7zVPbaQRpFnAvQ3O2UOtg/dqQPzVqN4yyOiuSx1I+1SCTxkwHmTPUGhoQ
G9XmJLx+O0kd6Xwj3+ElPe032ShlVrnAqoMiv0S0/ZbnKZ2IASxaFtppapVT2UmUxn5b6Hl59lSw
MkpaorQVQk/vP+RsIx6HumKqwfLg6KHaFHoFrO+cQv+i01F3mIqqXmxPKHX/w3m2/XkJJMI/Atoz
Yt09Z2SMMXh+S1zukkks8JqGiJ3amMtMqiaXjx2SKzPOkAPjy8xMJ7qkQW712dXDgj6WWUh8qJqJ
sTle3yy44tfaRkgaz1eThctfii7OjjFJO6bZzt+UbyCnf+lpshzP06mJcwy4aPzQTvokTmqx3U2m
8j+HDnSvgXLsn7aZ8Kw1gZirTbhvH//AZQepmueUi+dPCZqPIgMOdtpt5iwjwG8kHcWTi9YbHSvE
SsWDcyuk5Z9xugvH3ElpjUSvoMtzhfPXNYVoqm1DHes1o8OaQQhUg4vzTEYD4rg+7oUSz+2rh4lQ
AIaI7H9KaiVdKAQ2mjpeawl+Yxg6Er4xY34yXUVi1npGbmkiIplzX8yoOKlp91mI5BRfJEAm2l5w
48J2djo5EBuBDprWjfzBTQdDuvrQ1utBBkG3b8Qv9i6CIPLiy0/1bfNQQ6x/OTUIfsxibJCi8LG3
jvL1uALBeChSX+UsujHS+gU4mjl+3kq9Nwj7HOVe2YVrMjzwi5TxugsNU7buX2yxrpsN10ZWIXTP
l+Z6i7aga5reHqoYvyi7Yz2wtcjDHwWxd1mTHvbjh5UsCNaWulHrCVaya3AfzcLCSRwajh1nB4C8
EduiqI4uosznIz1md7rXRipTCgVL9lQIi3djU4TUt3bd2DbQBAdT4VPtcL2fUMOWeYgjEYvoMCgB
rbTQ+apCky0E21JqsPzX5slPlXC9liklO/D/baIa5hxVQYG9qe1oW2MQckRp9zDmksmmeImryOQM
y9nEiDMQiw/rZ5VUBwlM0T0J9LrAoPr9rZ0X0Nv+pUBfpLfZjqxn/ufJbIVgkk+8J3yNyWOYZmHN
fvIFl+ExOERcJYkHOtAX/g03KstO2irT/z3LUoQU6o8UySNeA5yKTaDKsVmGL0xBnoElCbDxeBus
+n3Dm10YwdTGSiGJRRJgDJofW75JvtpCm+9kIE5eAtv/LjqOXfIy5mq2T51WTfn+eYPkhzQQII55
zYxD7fP0dNeVor6Y9yNYaOysMUvCQcNnW2w5yoha54/qAX9FY6NTspGexSDcFFKh0Tx0MHVNCg8w
wvTvqKVFhfuPtlAMd1yKDytaT1N4xR8RLKi93qqT6mk3dWIL1HMhVnJl5/DuK/mnSV5N2COH1YWO
DlxkcmaH17QdXpVHjVgEGapNTcx4cnt382whP+5iG6jhs5ZekOXx07wkSgloLSyVzHwiM4dWXLOV
iG6tQRjmbavOvcbhrHHiZpcMzNW1w7KJrAsmxjWSXkgA6mOML9Q6dtTPH5gNjPQZMHFIWI3b9kSE
T3SojVNUl4MkooJ8qO8GCPNuZtRTXCOMgt2m5ktNBMB4nzNQDhmKpx/X5LGVygorOynpozSTmDHC
b7EVBYjEs1I2rwtKWLyzEMleboxcmaiWG/U7ZT63Kl2+Q5n2cjy8j9RpTu3vXUdCX28KZgwNMWId
63i0NF71n5iJ/xTG6SyV4ziUcPU7txsHjddag5WvcV3U0LTCmxKe+hfDzYAYSAfOFIkKzKMkVqSL
y8GgUzpEJpNZif4zfivYW9XHdCKhxDyLCj2izsMJ1FHTuLVaKSqGtL2PlLVvZDnDToNNW9gmuFk+
XzLcJlrWRGBp+okkvqL0QdGPJpcg2HECxF9HIQOteVFqKqs/EgLgxa6V+Gz/8HVZ1qv9sG15REM8
gDHVighEfQ5Ci3gg9V78C0SbE1QFHUYrCsLbDzN8HDxyqGW/5Zj72aaO3eIutgqc13Yo8+lw3Ksb
QPvIBN+WEOOSxa2SlbZAQK+RMg45p6jjfcXjXmbhIO+yK1vz0dIwfspfER/dyoGuiWruykn5WXbA
XkfR9k+mTdZkavf3gL09/lr7iQpZenMsuPjTjWjeUhBu3KvGIphiUcX+qn9Ufuz4FUz8k04OlmjF
FWYh16j3xnnTlIqtxBqSl1bki9oknXmjVs2S00Jx8b7Z1+bkkyUvQpXaQl2j0tk727aj6cIKmuMA
iE3oeUDELfIFknKAN1qLFnx6J39C7fFpqQdvqF6RIjW7m0YwoiUx/5Vk55DTAkfTwk/6eICNZ9b1
PYwon0In66cS5L9zqNQXWG/5eE8XOy4dSO2jab8miOB6K/gYX7rBc0ifGtehG5iPy8ntxlLPrfgR
vuJS9dSZKapERXBIP6F8GCnnynTnl5vGpewfstWJXfHYqJKFVjZV1JTwnj1W7+IHHv12k3t3vhaZ
UNJduqrOBadCdAxKs804bitr4Yx9K7QIEUklTfRg+e1RfydnrNOBBnv7ymBr4Pd67pfU7kpXbbu2
FtrDuADfWoXqe216Hgf442Rv9vrM5DlPBR6+QW4U1fe41XOnNUrFnFIb0fIMXs7M9enHfDSxnCYs
lPgWNLFRznrHkotIW7+UqtJ4hvi3zai9pA3HrG4B6Z/Ua4iOQv124R5867OHdQ4Xjg+m+LBtYSCp
M7Lv6DjnIpVjpjCnnkXce0xWAzRWyZspb8LRVd9G1fLhJ+hjISah+4PLWKeT8IMFIW8NUwLOtz6o
n/nbLHHKMNOZcmJRmhgo6/TDoPICqdNnSov5UclQCsTr5EE4SOGpFbdMy4t786e9/heovDABfBLf
p4dCr7g+EHRiVxMyUNwzPcpy7pn6OuFhYrz6R0qufBdBuwYWJZL26dH2mKzVcurvPSba1KYjO4Dp
KMks5ngrXRJyGb6uyEihw3z1KcZjvqhV6K+q10ak97mPc1a1ixceAjK15QOKhm7HWr9Yp9V2KkOI
UhS4/oyjoEKrpzoprOWS46eZJfbDB/PIUGFftzGlKEkdFDnHXjK0itlnPgfX7VjE5FLyaxH01xAx
1T1MuyApnKXtzRmppdpjBZMSSZ63xvLocTCP1T5/uey/sZjxML05n+jyTZnTkrcvLP7UsIAhXerh
U3/WJSWwmyysfvC7sIvfRb7/Mgmu8pO/0o9CB3CVbgGWe/Ze7CIFhRRJ/XPi6KEx+FOm/yUY0HN0
bbZRycrJ80990xxHKe2Ns6XoG9HRZgEMtx6OrzI/RuSWbFkmsJoCHlpC5mIUNbgCQeM3J1clWEFm
0A8sSMiwNSotHf62C+BNzO72S58Vh0dKwGsjZ/W8VU3xb8Hkqn4ioooo8857Tq+HxVM5+ps16gNM
Tsydh97JQn3AFhS5eiQ6vINDdRhVscFonXmEE7FI7GnZpzfV+HgvRxrv/KjCdzEepM7LAybyiWHj
NrJL2Q/QCITk4AU5NWnInhISbrqvaZt+O6k6qiOTFofzuVIYF2ZJVO1ZC0eTOSZwkjN2iDRLLTYZ
VZGropCpVyaUGYO54PQw3F9T7bR4zhVvUyxWJNlINBpPO1MiG6ntZCwwmjaZbGWg00KRx9LCKLfJ
qJgKj56rpqvhSSBweeFt+Uv3UCC4iTpkdXp44MraXlYgPs88IU54qk3TxcOV8zgDQk4TwFa3xImT
OCpLKiNOex5Ix0nFw9mOBQPJM/7Mdz14kVZo4f/bF1p5a97nKXjvA1sJRbX7qTdGJjsZEL0T9DXM
zjG5BHYZm+wkt24kE8oN5/TxhTPoN9YUN9v2X0Nlq3+g47vZeEVtO3MosJjc45QKcpSiGFXJHE4T
3SNByEFYbcbQwv2RbdCBSHZBsm0X/MSTmoeEO/FCGKSLZiFh0GnmTNkotCkkRnFT5riip9Hr3EvH
j+nqg4XsdkVEMtmRmTPAsWyi+iCdYJrHtzlwJMohxBo88icxaV+l4b+ZZbl2n09WOdBMGlLwWHj8
3Ubrp1wbCXzknaFvo7u7K+eXVR0QOQVWCCSZUMBaZ0qe+COmpuoGCVDb4FlgIIcU6ksyYSPoCayq
tq9PTsK/hNo6NZgodDXb9tRdksfNova670h1hKURtvHWPK6dWU0D/BiUCx6UWua/O5rafDO3N6Co
XmV1vsUJcK4DjYDFl7iPioD4YhSELqUZzB7vnzNccOzOtu4NI9zERF0zm8i1F6RwMraI5Jspn9Md
svk7pxcKM+Xeiv4M3od06nB3f49ckmpzN/rvwkecX6mClq0M6EFsb+gS+R+b8OlJrGAfIccmpYmw
xI+ye9b4LwmYCwvLS9q3XfTGkgA6lp5UYPlknUOMeFYxAfwt2Qhiue7a7Ri4GzmnnUMKNZ+bVfK5
GIDZo8T73fuhDzrdvdBnfZ1hNRM7Jqeiv8MV59rRyY7BLYVrDjNbcwm6rUF/erC5veMrcsZYsA1C
6s6jMdeKdnVYCAGyZAhrBpnpCzI9KJucrq4tIdp/cuo82pE2Kn/B4cL/ErGQu2x59aEPWidv16Q9
PuK9plvDGmI1biRRQo6FQYwx1STXuUHRMDTFVMe4poClATOw53Pj/Laz6d+almETsBMeoRBcbKyT
9bgAOXhv+mbFtwInIlgn7he9S96uoLWe/FuaGtjxvEkbo66M1DZ+72RA0z81ZDZfZAlxpHyGD+Uh
dp74tjf7q1SKFw240kcRnGMS1Q5jqgW3QKvgLSfo05yFbAE90euOlv6zHYnGGHPmqTzeJrt1ZOM/
vkJt+P9lGJlVvvsvCuLAs1Nx0gNE7Iq4a9p4U+oQgUgVmV5JpJT8PcF4o2wq705utHcsfQ2SBef2
wP2w8iDAEikxx7R8NzTLMo4DG3Az9ntUVNPJnxoJQBIRO+IIwsd86LkEiBv1MtOJ2CPKfFc2c/3F
rqNds4lMoB8JNJqmuVS20SYS9ytVxa1PGEiPyBP2tIrQKZiy4YuLFu2vIXKO7arEBooMIxcpOW5u
cq+QMLiLxwi8e2QTM2ais7UJ6VwjCz3usnxj64zpNVQRJLAgEh+SzUkOCD6B9rVJGIcc9zPNDgJD
LobK/L4paUDKm/tpBq7GQNpevGD1sjcVhyuNkA3IDy5iu2V3593fQvJsugumJTPwdf0hcHWf6btq
/h6VgJmZ9o5yhC6z5X4m2SrWLMOsnSGV8LfZP/nX3jmqz11Kwi20SKwTLFw1CUyO6AXXnewEoCM/
Fz8LxeaT6yzDbvpiF48DpObvkb1lJ/1dF+eqByzILoOptuVZhbTDF2W2zzLtjS/QV7RPON0jAb4T
3QwPQVT1dB5Mxtc9FPXw+qarRCtaZmbhdz2BVvWNFONzw5EFW0o5+qP7wGeuVk0VdjDpZAtr2ksy
Q2MwsZeD4hjYcD5SYM/armAQxDl8d4oFejUuQyffD6QRqfKS/oNqIbY7334W2GXBxm8TPskBU1Vh
8uIVXo0Tfi6gpc+fLeaV4JBLTL9y8riEtHc9tVKKA38objwbk8Wm7C/0n1hhleTBa6lLO6oC3Ie0
NO4X3UhpSqNr0UnCfoU/oOjSrceu7EjQ1wKzrEKMi91+ioR6ze2SN4C7L7/wep+/6ffUhig7VAAn
eLdEoK04o8tUVMr392kRPMZLwlTIQ63tvdGw3n2QQWn5OdbV5WrIcpZHpHc44wNusQ6LzAUSB8YJ
g02/w5EWC5g5EVlzSq/Ay78cBduCJ79rVslRJSHtinMOIVUuTrsGk7C47Xppmf5s9ikGMFfA2xIX
bZI0jHW7ec/j3Nn320RQTYd2TnbaJjISMg5Zegj+dfOWk4yXdS2OiKCSyFqLcaBFwvsTJ3LLAzSi
76vdy0knM66vEHnCIju+oKX026fu05XMKNzmmRJo0caNI1/pMklb7mRwN92ApnfYEvTg70LJ6HrC
cT15vZXPe0i866qSh9W06e0RyJzn2SFwpmxnw+/19c2Gld/alAcrZbo1Zn+mxzHCrv7uNOpOLeXU
sNojlsTNFj6iIB2foehGLFt+nRSvk74jxZLBl2QH0Hd+WU1vfUuT2Ntmr42E1H6ZjEB9vX/ja3X0
ii5+XFHSMn9x++4XKamk0tt+hy6x54G6B0rcbI162q3GefxQTXAUebXm6IVH9DBzNIzQdpU5nq0V
gCUwSE2Ko/HGDgwe7/EucYgl/Gptka6qlBlCe5HxlCs+wp+Q+SM+RLWcnxYzZzKHrUQBiKIfXqEz
amTcVXgNmboOy7ADk22YFr9Iq+I9KOCECS3MTzor2Gpm7FCwvYwuN8MRnB9JpsG0QJzjvZGxkS43
LMXWxFGH5X+oiTfN1D1zl9AQ0p3UKxVxozRxE+P4dI30wlupsA1Ywxpn/JE1JMV4yceTOCYFphkg
gE8hnJiL+lL3wMbGhbft1MZ54tynohTgkyj/sxxmHvxxg5pIXqmEBN3ggdIrV27v5Au/jdzsQaIZ
90FOUpiVRttb6WoBJaf1XzUcnepmVXlhbI5uXqrrfhvqd7aUExXGZfthM63OKAFILa1wxuZKrpgb
4l9qVuT2Vqc6OF3lzOZpjmS54XwFdwfPa0wYngnWCW18U3XInF9RSTtTx58l/AHDXubiO0Wy2efa
gQZDPmJ4cSA5lgSEDvwFREuq+aCTGwCrSonrCdZqZ9VnHNMa77vbfoadiJRHZ2Z5/zWbQ2XUq4aG
xpgjG2fTy1pmiTTQPBEt76bVEo5Te7xlThyA/VRbnucBOMPN4El5wRmyJUkE0xTBIOJUJHyH+Yi9
A+ZNABCD84haGRMoS6Z/dtpbW8c6BU1ehWhwNAu7IXjnkaEGlt25+X0OPgYE9CIxHFOo46Ak/DdU
T+ZWZRRMTzUcp9naG4im+9b1Usofqru5htJDhwJuPIavoMD/kFQLbRWQL6xnm2uMAQjf6ESOw1vJ
o8x68zpRrZUX1PMw5R9WoyAN48PJVCsWxS9gqR8n64H91F7dVT4EFwCvXspHmDzKejWqoKOzY1F7
dnODT29MGhbqKRIe8qTr21u81cug3XR+cTtfBmj2M73HZEgnL8W8mEFP+LgB3gJLhhhpmQyqcJcI
PgNcoKntRSPjr8wDrctuaPrDx0rY+KdwoAa8bvHjAvoAT/VP5P3MBIaUAAPeNn11i2qgbUoLsTrK
oBtEKvwaQXLacFj03j51XRhavasAAfsTBKsXJ+Y9RIf9ZsEqdzuiqE/SButGvDO/oG8dy6S9+8Dk
v+o4Tr3RycGPATD/vmbYXY5Zp7kQkgUxsUniJR+9F34jQU6pvew4P2gOT+3OswQ2Yw7y7jVf+28q
c9REcyiZMcPkKm/qiIBbrfiYJvxVUzEWXq9ctwScBrkp+h9AupLuJLzOdUQCHk7Xw7SouVcP60+m
BSGns7+QYX1rY8gC71IsVn/8ryFKOjeAf1pekE5jyFjuW9n4qCEKbPVlJ+16+2J2HE0K+m9Uz6YX
5Ixf7epDSWjkO4AHO6CMVE6gs0WUr2OeYrUHnLU/9Yz947238iO8n/1Zsu02dr5uMwZEES1YSKY2
MNM3AJKL+nSvkTmdiq+ZEbT+0etshLnPM+4v0ItLqjr8/orhBs/ytoob9OHBYnALOEWBknYRH5kU
Sd8THhDtfKH+JJ9uXnQMsPsBdWMAAWEqinR5NUg24Lxj/OuKCvc875NLUtCLM4rYSNQsMJGdEKTd
uTnGwgTsuu+Mxhx/sAu4y462Q7csvcjdfbq6Q1atkZQSuGPqOYBtNz3S7Ch/AQ9WtRAG47Lb4MjK
6gp9nPqm8Iydmb/eoU7BF+JQg9FA7P0ersKiMxGZWUOpI249T2Jq087w5MmyYwm8XwYmT4Gqeazj
hejESGIVDZfkqlmAnNh0mjwLBBQQjXn3qwnJ60InPViMF+SNz94oW4yXufmQZp+c6q8yaVbBjgwK
vGxFt5lbHWRRmesUCSPFVYOWSkvoEoD3cmtxacy5ZD73s211C+kFTnYXqRvvtWfUnyk/oX7CXOQ4
ZxuWTazt75GSujKtBJI3pmR5x6GJgPmINerrJMe2WTvt21fyOvu7shekNRtsHvu75QVNJEfdVx8P
3zfEdvM+Jdi1fVDKtRVCpOrb6dQ2eZYxk6wi3w7F/4liVI52mRevExnz5umsT5b7TfP3GJlNYiEi
2Hwwz5ARA86yjkzUJ1Nlwu8Mk9YrxRcmXN4juTHUHiV4WKar5E5CPqBJO+49mbFP0q7k1L0acB3A
U0E+IjUL0H9CbM1/Zq9tCKBCaqhNq1CrlIKUPT6VzcYiOKMwB7/sbfsNkJ1pOH6ID0zY1JdX6pCq
SXSojnQqHfd9owcUCwMToLmPwH29a4XLOQLijZf0J4xkD16F2CJeuBOVWGHMVuk6j31yMyuxknEj
8yQ8KMhmN4emCBokPccxSOanPhTtLSn34datAulxlrVgPhilNkVMzJXTbvcJs08DSY6imlxe2XuN
p4Hp18WmHNFBOnEjBmTAA44AnQP9CsxqcBCWYH1Xa2MwY9fX3Td9qgwv5FztTdIQgRIftmIuVrgZ
LmiFZRSI4twuCXFhFkJG9fYrLIz9gPA9F+6S7dW3EPN1xQUnsGtkgq2vpL0AynFX0qaVPrD8h47n
WpZ+3odEwSG1s5QjAjTiLec+bVF0qx9LdpVRjoIX1U2dM/SVe79f2d13bwj+tyyd3zBKL/Pw6mhv
KnBgnswFEJJ3eJZUH8pH2/RAnCE72SVlMYn2mHVNtKaODCq2pjK7j7y2RZQxKZf+gKTsJB/2RHTW
gHyS30zJ0YYtUkvVKigHIGzJ8tqNfjtFk2qg5Hz0UsizAkqDEIczeoGyAY4t7yt1mNxrJgjKpjO6
7lOtWidyCcowKSZrg6L3wGOU+ZlkSiiDdht47eHxfki623jUFnvoKwkqo++whNyrdZdPmKrrq46E
Mgy/tbbh0tOHnzqsqc9dY5cadtybjInBjkprSOahmzovCi1r9FpuvDUdJSGeY0ZuNkhWC97xRNCI
X6Gj5YXao3rwTBanIsS08m8CE+H2UMQIALqd0BqXtkfthNvoCEr1SoUpDj1Qjh5sVfdSbRq6Y4MT
peVCHYg9Yjj7OiOw7L1A6JXCgbsZSdsiNFgh1roNTFa9kfTZV/97zEc7XetUSi78xQW8utfltXd0
/r/DTxwpZzwabOD0dQJbU31fULt4Jg5ll45nCXjSj6h8htc5gUPDNh787lanpVw7+YigF/eTk4ar
X5vtHPxuK0fFxXRCcum/q1PYmVnkEFMBT/6KTaMYM1YFtFUEk4pLZSGxTtTHHNj/gH5frD/JE/zJ
AHpC2olzViJ+NtnlvRhr5/nnWdNtp6HDZrA1um5Bvx1lAZVsx7kExhc03PBWbEi96AiOpy1C8FB8
Tb47844BIDDHXegwG+9EJLnD9hMy3xnkz4dLrGfyI+OgJMfhlGAYl2pvgmob//2Y4uqmn5gCvP+b
4bRpN/K6ZHFBjJaNdGmvimO6WsW8Oz/c7wH6z9Nc+xtT3KtW7wjf3GUxc7ipVxPP5y0HTttXATJ4
2549iLaMqPAs9EyX1TmR8e0qsh7TPqMVHVQEoyEwQ/CwLgyqldwLebKEBqiLwzB+X2pM4MEuI/rO
nalGyYPXX4n6Yr+eoHxj27KN+6ajkPLDE+PJp25IYiMar+Xq+uC1QbUSyDHzYrkBOz+BgEE8rtIf
bqUEAT0+N+mNuGA03ax5HFZ/bKbT1/CYLhWW8Q07YbnUpx+0hfSfEiOWOuCLN2L5J8p/NPR2zmqe
Myy99N5Q0LrgsRRAQRlCZcK2AReRE5JiZVlwmWm0y1gPJkanpGb0MbQrtcqzLIlkQ4IiHks91LIO
rAHXCB6tPQ/tjd01epi/uI5w5GcUcCHb3vZy0lqQGVWCrzAGcVtnBN0MVBmFruaMBxCMN5fVRv6o
zHrFWr2g+ISOrEU/0HmJPQdM6Vtj19BfIeS1BlzHbWTEMC992mHYmNOlXB1HA7hTp37j7sCappub
Mn4+pxfSsVVeIeyKS5nqs4nvaqESqNy4Gt89rQKz5nR+i1xAMz7BtVAxahbzr1p3Yye0CRzCK6OB
5BQdHkBD5hCr+K2cRbmVTNz9/1MR3XvQAg//HsLAa9JR+nW3HVfzQjLF9AItdDmmgJPjoJkhVW3t
Whcr0rPgNsTF+P56DTyAWW50753nmLtcJj2k7U4orJAmKR6NQNtEesf5X53ivmRmlLEvstBgQXg3
W9uZsiEDEav9u2H9bFTfHjA8NOJ0o30XvqWXjAn2ghyHQl0ARmy1wbWp0+f3FS+HlvYv925UwvM7
MMqSTMPX8WshjDvMsKN6QZiOTcZdfntLgzMGTrzW1Tmt1OoAnIwp6thhaj1cKwd/272mfbtOCzJU
NUIPi4np60bO3eIbbKfsbVGM+I/oORyRXV2NSnWhRx4sZsUULT/np7G0lLDOnP8RYhJKv6YKKO9L
ie7CZS8KKzxO5FmyeXNOojWdNcbRPLoU95cjE79/Og4gwUt+H9q9odkNkNStvZO/8wHqceKrJ4gQ
1xmq3qw7nWwx1mcFYrRu1LIFoAoAbyGROzrIbwKr2aDQj2HvowvVpwaYApy2cB+AHU2MU0uNd9T8
XrNAjfUnkD0nxtn31vBLlRE0TrVD7EZkTjMnPDFQ2OXqoAMdLst25prdYW8afTe8qDZ9INwvysEq
ki9fR8qoXtk6VEKapqZcpYR5QhYz4pu7oP5uiWasy2foAKUYEOCXXupQFEOX6QXPqqR96Aanofu6
Ht6LSY+yrlLJIu4cnuiY2NQLtsWX589G2FSwag34pZ55BkcWwnpQP5w9OX2p/FLDU+QqxORnA44S
GiAERAG9g6ujHFfMiSfi4KLd5x5cDnHPbeK58go39m3Yi/00tRhRqMpIQzplilUCv7pNcO9H1KW+
COZMHKHEeYYyPl616ZQ/Ze4mBdIKFZ9SAeIDBdfhOo++kpamuhwuX0F+zrJLrvyJKanpcChyyVQe
m0o3R3lkpYD06iNu6WpYV51dvu6JlNaCblI1XBfoV16v4/Aa+eQlKb0bhZTK8iH36rSc9Wq14xtY
kKF32DoXhe7rDmCrQGmdXK2C+98Q3BcXsviX+fj9cK5AkNYWj2IBC82bZeiLYsHEElxhKzVEbkb6
HS6iSSwjlg7t2KqU33p9RDqG/nC2Ymm2PYyz5gjE0XBsOZHrVCf1RjGCxfdF7OLEwpPVgta0kvZa
Vq82HILj+63HUbBjv0jx37GWDOf+ft3fy9uKR7Ek+PQiVVaxWSaFaANSEEvy4uVcc69WEPcQDH9Z
lB+NoY6Awd7soC8cuo8c5wOEREcKoJQB5fDfMtxlu1W6FkGAa4JfXBaNGDTxsBM0Vp8PPkfOSsSf
btbEe5CZy7Iug7ZAehz1v7wztD0KGGMPsXSxxExWmRJyGuVq0IIdwi7fhnPQsc1unGWFhvKgLRFq
kigEzfKDpXj4hGj91T97YaXAKoacyJa33bJRqM71x5LpgnRSxmN6ClRnI/J38XZp+sy35mBHxhJi
HBwceNrCYJDP7vY7Y0K6y5H0PD+iAKTpeJD5Iu0Cb3ZB2UtwgT+lLiqDLNVhSOxGHj/8BvXPDZWU
QGTopmv3EkqB4LVwCZnCDhcmNliddRPnDNwm/43MBnWLdFnfKcavGq3mLKPVtGW45/6HHWXVWauh
xZ4Z+P/U8pidKBodTVV9U/vWin11xumU+KQay4CeDpypqylRgcXBcuVWTm2WoiXlc6rA8pyHQjzU
bAV1KVuA6/0fyFtioxSQRvhIIEArf3JR/lSz7cHQVX5ybs1+iiBXCE4xogcC5q9CuJO/tovbY+gV
ZF29wK1dNijlOm8PJQaf2hybT/TCPu+XdPg3IM9eRBnYnzHtoILBUANvBlv3nyp5dM5ltN93wa+d
b55tCFdqcsA7d3W4xpefkHdFTIZUVMC5sOhpWWnvEMTmo7GzeaqEux8v+c43wFZLOEyh2vx4XHNy
R1DcZt0naKYDzHgfS+cQ6H8UhClvWDplaawWllkqe7gkIv+opgWvVG3+VTls4sdHaaadufHOCH3f
2MHVmoIWwjuHShx0vylUkCdXYPmA+Vi6xq7bgkOkPLUcwrfH2lLoc8TkO8PhsiRVRXZWu2AjZtkU
mZOsVXN3pQGlDcszIPGR8S5FxFkcI3V6hlHCa8Itt2xvxn4K8Oo0VaGI75QBLb+9hH5Y2d5OgW3I
onNS4Kdx+n34SHU3zD6YF9qKGRlrqlyb/BUqchulKADvkdVcQxlBTSsjOh6ptXC3uCSerowLc6Z4
Q5QITRDWx4DLhiLyO2AkS2bZtK7iEMNuSlyMM5SF8YmtVECSv1FWwKUieDPY/EG5GEZZbWWdbkOL
vqmSbFWXCEHYuu8BfNHfxfw21IvMLELOfaHDXxyZp63+EJf+HtZODr/PiBSBkjkGctHsGzEogli0
F/LhZ3IDdJJ0sO+RcZSJzMU3c7e8FK+XGdXcv/J5B37/wo2Kt4ArDT9mZJlkgaL4udwjLbld2qg8
Xx5c5b1LQ7fB8DwRsP3cwBOAxzDNB6pZpGRedxUUY/e8lLuvNR76IqzdvpG72ZA21ZqiERyPs80Y
E/o5/W7ynMCHZ53V/Abq93vRc9Mcs+cmZyJqE7UAO86RsGOEJoYKxj40z0g8c7Iox+EDQuXvf/Lr
rdaope+TB8H5b/okEvKzA7c80+EsIs7pPLor400qTJKCEJL58FVrD7gKiqq89V1CmvhV2X86nLPB
S63maQ2Nu/snQDOd/wtbGA8LE/IWXWSeyPlAvJmK1So5CbtIdC6gqOLng+0f73kBiOfwiAJltV+q
5T/aB2z7Jl/ja6NKldt2nElCkYAeIxDMZ3Uzo6a65PBZ7j85MKn3oqSX72Ve7vE6IWJaG7Idt0VO
3aizyPST7zq54Ht5d4LZjUCp8Rix4wYD+f2+dj7c8XJaQEm/sGIa2X3EUTd25Az6ZG5BfN6WlxKF
4SGa8K33SBA55JO1Eo30wyq3WFwxgC/vuwnH66f+4JWzQt3QgvOkbuGbryvDXapFRay4e5YpMykI
T4aMeJYr/gF/fM9pE4SJYPznvUUoHOwm5PzcFQq8s15wYaHO15Sn5dZ9JVlNpVC/7gr4ydsKUfQq
4VbmFxzPXTKBCXyUlCFJS/7tNJjocn8Ue4ripFYuNkgdQZ5lA0BbE8Y7xE5Bm/P/J8+mwOemsdUd
BOv0JgJ902vhHAaEsaYT/wjYQkHz4rA5ixlN5kkkrCIsZqbhoGdV+vtyNPCuYs5au026OFNx5omR
oWReY275nzj9QEgkS6U/58l6daHRAETx8c7wIv8IUwvj7kuxrwnmpjGN6fYq2hPSX8OVo/PUQKDT
ZMjqR1RbvgoR9z2EsdH2p8Fvh7Fk8np6R0CeYM1cS9ThuRl2mXZyQEnThhSPHmnVZS+16YS//EEd
/exV5RJNxm4KR8RncIvMm4+g6v8gkzFznp9UEDexlURqpUXU2cbVANM/q3tzCB0PH4r3bNtfMihQ
TTn4M36f9qO6r+0p312TeF4MZcJIYG9BQ8Ic+cyp/xpC5fAmaEiYTXkAJDnn9zOAQ5aTCMFAuQ+s
m1h5zC5ynwa36o736CgYBkvB5JG5S1QKprzBUAzwUk3koZqqUhoqE+MqounVkCz9ZHQduJ89XZo/
EYDmglfbKYZwa1uwrc+Ep8nPWw+43NjP6vXvDoN6ZtsXYN/+dtN3GKpYAJsu+micGQHYn8WDJ8U6
NAuc/Yh87+BeNFlzZtaIZN8txDnpmrZP2wfVHRnT83njpGW/dl6K9jqn9vSTnpLC3MrLyQ6yYHfN
wa/YeVFnTcdloVFYO/fU9UQJsvznSZfUyfb5gB+Gi0JK+ApbVC4J8VE+UJFLz75qtVjQw7b7kT6x
CfLI0+zJnH+Mgx6rHcYnlyLAqu1fI3RyIIlhnP9aHtYm+zV7ch3TufnoB9meYLYOxMKKAlVug4L6
4gQ07MCQ1xR6uJCZvzKy8YSDnWwAYNU74zM2jMHh9exJISf+8IW4sHx1t8t1ZaUrIlqfZu3KsVeJ
9yLR0Yy/+mp6I+i88HgjnRAK0swXBQJBjvEqFGJ0PU3NV2/DwyXZxgYvz3VN79qPXxJeGrfa/qW3
fc4HnaDN/1kF9i6OnW00Wc2rYlomMicLl0cakNQqUptfAh5/mljBj6ihWFh5YlIcqe4lB4KQtsnf
VlNmXQVMzmZExYl++0XU5q7o7WcK1KObLWQGAzbKeocbL1gHLShlNig0Qz+vIrGALcDXw2MsEDTL
milCHIL7FhLOI3tB1hiRuTh9P2YDdz+lvw11IzOL5exdaxTmpqX8f8RiM0fhZccayDWOuMXN1+zc
GqLW8coZbXe3pawowlQ76z9WVkWBYyPv3KsI7OQj3rtTPCVonKLlj7L/rUMHHR7tP3IeyANQPi+R
QtcFDMBlNZDX0GlKM0LtC0sQrnH8MAY83pbuTVjxuangZ4qnyKAsb3utqQS4k3qbdupCALU5fkbG
biTKK5+G4H/m0tmVqo83qs/qxTcrZAzI3xZ8xzXWV/E+RZONGOrThcSskomZKtmh9Q5zAflc5tYG
hUX8lr7UlViP768Ljk81PElEpl0ZFxJq9DaIVEADMkTR3PDKKloNrPUaq8H+eOpjI6rsBOujqGQE
zKdXr9/oHGf0tA3X5ndDa5++DVPPJDiZS+geAGBJEkC7P4KnHwiHSxtsOyfE8XZ7hHZaKHV1pTuW
7/e6Cc8RImCfYPABhEjdRHFofucMTM8HAYoZYUweUGpBxZEEp1Jcgd9CM9R8AsFO6Wr8fE282qGY
vUkQ6rdxeJyuqVcn4qU88fGFSU6bLWtHeEsXl2rKI4bsrvEY37i82rYaj85gp5f3ISpq2QnOELMV
ujpeK+a3YZsFh12p7QL7aKjgyB9H6bY17Dcd/umpYEGL4AtcMrLoRkxoG7J3St1JfeBrn1lzGbQ3
3sP9sTHpjlstV1d4mRFwAtXuyUmvBCbSxIBt58exixjK+HmGaNtxXzIPgLuALuZeP+SnIVOH5/3c
OGP7Ujk6gK8T4x0jVqzvGIjvGLc6AOuwbjRD1W9w5vaxtR/XwVIbsSIohLlIdcx1dRlVurznrC5s
mAbWMEcHODLZ0DaZbMXiQKX7vIAVhTz8IMJ/awY7uLob/2CE0WXAUkH5FsvtQzFNejihq+jPLi7v
NF30Gu9WK+4OPOy3Gk4+pm7PtUGxas5g9mEQF7BZ5T0OXs3KGNr4+RK9gLV6lfwwxR/E0eGu6NP6
w+tyxziG3bDuVCLzgtKfbxMZRD8DM11ywev/8hQgfH+mbq2fuSZIgyCdpzW4L8BX4ODRPAsSVMzm
nmk6PMmYIeOHR4jKlxtrmukDui80DQt5ZoeLDBfdJ5algfjdx/jDtdultcuJFELi8qAZPhuYRryw
D4ZqAKzRXCsRvV7g0vIBmEEcDlj+2O6lu+VSqm3U4CC8I2dD+2EW/2Z9RJXAEiSsovJ3HXchzCyx
k9igLsX6MgEDUohH5KrKYAVE86kTA8RduhkpzCWr+4nm34G1H+LGd4rycSkbmKaiBnn6n3RJMR7v
miWz5cUJnJtbYWiF9eiKkYNgSeG94IdigtWjUesdBzySQJ71d5MZj+lXqV4Qi30UdpLpalBW/YrF
AJqeGPB0QlfXVFaf+P35+HXX3L3ndApXp+AeOQgceTOImzD5A9QzcbueaJQpL7IzW1vZtqwLZGBi
fcSJ+vQ5VUopuBHU4HEciUmgKiqCNAlTa6lTnJsBcfOGU7P2H5Q/WSsXFjXjVja/OUxX8dUihG5+
2+yIaz971+Iiz6vuI0A9jcEQYCOEs+essRJkdUxNhzGwaO61OyaFgjlDGlPZ1W0VTuFG7HtuC3q0
euU1XQnT+0enqJ+p6KVXmfgrrvsr26Wme/3BJBUkMRl0Hb2xuiKbCxcb8fFgRHwsGh2iiAJkoYFo
v1uIRf32Gql95ssUGqFZ/WwFIH5nug6KonZIdVkgjJoPbt6H+V/ihDIOAyO/QaHWgXjqLc9aNful
pdQQDHLQuJQzZxh7qUjHCddSwdvsrgeIF8umPC0JgppoQ/evHbnLAgumu/vBiLpafL/sJdrhYbVq
revZzrkCiKyFeiOaj8APsIl/KN/wzsDYc+H2gMZg5rRAa8hRJ63UzrLr7mYNg3elz5q3APSHrTxj
z2AnAi5+IXBr76FF659QXBpeQCfq0mT0CT9bnoJidCo/A1BwJf5o7Vuj//pj0sS8UcvUOxinln+s
wNm6YQDbD9buyCtUpqzhh9N8i5KGK/mJOHlKaCnP9zePNKtBxJdm0Hb15qEIBD/Yji3cSPaXUoco
5O5lAv9FVf+Cx0efnIKeu5Xmn6ONEt0elM376/TwFfQHgzXr9RgQF47QnVfOb+e3Ohu8QWHsyhI0
acnsl+aIK8rMNcbVeeMIosoXqWWBwDIgrkZdbqOrOX8sZM6oyLBR2n4MKu46gmGY5rLKNgEGgLMm
6I6pml4tCcIQA1lJhx9HaIdY9pyDJUsrWCQmclgtTgxw8qa6p5D4CD9ld8Ghy2pGWsNxug5dUdxs
MWbbMUBimKFByojNGNx8ETRauwfYNUwMRhJqcf9acfA51UUhzC5VT0iv3YlZp4zLNbAh+DZBVpUC
1hW3UwloE2IhB8TtXTJ/IVkYD5/89mX6PrJGyiemcvmbjaJLCSOvJavEsy22D71EsXdWcmuJ29Xv
jfIj6nckRKyAAJ/3GCCEeT6HRc05uVoR2R4kKr5NGMOjpP7Be56D8M+iDuLMxJi41ALJgQ+y6Be8
LGylfbgRU3vi7eUCYhkVC5XuMic3evlIJzceKKspnyByU+c9f8Z8qgC7ys/ZGEcNC+iRznOBujnQ
UoGTv2yqPELiD5bqC92qraKkpst5w+jzRQ14y9kNJTHrIqcFGsSp86u1Fs7A3xQZ2+qwxIA55fZz
lHSKeHiW+hgsc3dEPhSVeqIw7Kp35Dex/AF3YmcCJBbuSqNjluwzUNIdNAhFILsPIj83geauCdfT
hika1xuLEv2JcL3mThJglUy9AZIyfKovFGEDdYM+TR+ikApwez8wMmR6uJ5y3zTsA1HQpBN1/fTU
07in6iadWqa3+ug6X4dm1Tvc/nraU1Zs5uK2ruBWya/eLXuxuNf+oz97nyqQMoxV7pakRSrnDra9
Iy1wNYjPPmXyoeJL3Veya+Ay+6mEjODS17LcYvsxxS4bF010G/CKoEUc7Wq4th7HfZiRQH3rjtER
vJuU6QBZ7GOCUNuIk6Ca8XMQejpnfuuE7r3fLlhfTgWFhJVcb1kg48muhew3gp/8It4y8R0jZtte
K3poW0OGSEhgCyx5bP+xM39zToC4E2wk4yaKJjdzTQkfRlu+I19yGrfeHg/uAQ6fDngErKDjGdHk
iWPFjZiAOTj0coIrChvVQn2Oyf6W3ClQLe67dpuklqTOIL+IRJGHypX1gavafNLEpXVfLRAbzdhL
r7xEI+vJvj+glBv8uQKm/fuP4Fy7qgoVEgxUTCN1XHonTzhA/m1tWdYpKsDUbZLCvkgKJ6MPEPAt
VcH1X4N6r5e01TomyokrKQANlpdsKXKRCd9Cb+YZR566ZgcrfAOW0Ct4RMl8gLpcxgEf99YgDt81
sem56vESjckUoNz+aA55XhmI9vyMbiOHm3/HWu+ZI0noljRtxI08Acp4t/JoH6o5rhdEE3X4BOzn
bSj1qL0y5g22jASNOwnqH6CcJieQT2LtJfiSNXUSETcPNnH6NMZL/gZRfPGBRVY8DCtfgL8MwM+G
92c9DKeyWTZO6Bizm6OVv6NdWy63rSvN9sgLdLhJM0I//28X8dVLIi/a07q/2fiuOc32S6XQOdwi
eOLbC1KNO+i+e1CryUA/MsLtPRNA40q4KglDorPo6mhXEOgIvRG7dk/PnSu0DhbmwJsPQOrKgR4K
kyBPv4p8EtWxSHt9u5ZjQC17U4mssHxlbB9lq7Si+HY7JApu/Msbn39YI/KDegA6Dtk2S6tUzGjr
jrc8PLev9mFW6E4iiv1m0zLqNiqWrruee5UeUgy8DeqmA/QLrfS//+WNTLtpDVoUn5sueKtfVJOZ
S0qBZ28aql5YFr91RZk4aovK1iTlKt7dxUkZfLHHj2gK5wyzCu19sxaCtYrnI7qyeBNQviniXxnI
QY21usnNw7ZBSsdkdr7cWPtRAwk1S3bqn9cNUKQjagRL8YXNaP5MD2r9JhcU3dp+E4OEFbLSHEgk
Am3A3IQ7WS0vGm/GTGj2xE5eJCHkflN5pfJQzAwkAOoUuQjc5i0nfmHRT5VReIfqNDqQVKpFAuyl
JDiAzG2xmXD7+HFt6fqnmovXmWXHZGrx0oRaQcF9LJuu44YfH/5SjyfD0WpWvYiZneIGCj4/BCgb
2KsKnMYQRR4tkjvk56PaNso355NKZlETBui85QTPOqC/cXOYs8cz/t38V9Oq6L/bPc/NOEaVUIf8
XIMyZ8cLjjZB/eJRUQqjNjWGa9urDZ53xhHrAssrHkoqtzG7iEc5bpGBOa0TR58lHf/gwdUO1gjb
z+lXc3MZhXTrIrR175fBL4FElJwovLGXF9JzmjY4hGh+vW8EVEp1NmlgHDhhikWf546hizorntD5
3NRJqArcyN3A5LCdClh1xf2UvPFaHFcT5lMeAzS3gCsCSMiz/VGEJIuQOqQ1dF/9TkX3blDnqSdW
BgrC3HmMKnvmFJq5iD2sTE6KoXdqhJRkeuyXMoqdDzvhBBDLg8+ivc4tfmipqJzrQzmfpPU/9VVm
3SHFgDpNXvyZM2OOGgW5sw10GKwn3WVyULTctE4YOhi7uDnmFL48tvzaOnVsluuRahIMWyQNhTmu
Gq2aDlViVMKGEiqWbkOtNyv3L6HpM4g75UyFiX3AWsp/tQF5gg5jN0q1R9UH+5A2vfJ0iaEmKq/T
N+R1HMShOzad2bLDEAlQMlgfixEj+Eftyrs88sIhRte9R/Iya4yhIzA4e2aLP/MP6Hcp5hHlaUjy
tljiU5w7G6Hp/u7oQMSQHmmF0CWeKnU5GUbMvT7fqz/3i2AmCx5hjIxnsnXHVZ9ZVqFN+x+4ma6R
DXifLpY6dfHLGlMnW7GZd016AKBXxO81NNaakF+TwpqDvL4VgaDAgEdZYm3sqI63UdCLjYNpU6mf
KAvllNr7pUTghbuqDfN/W2owJrMHxsOxsrs0aiyhlIuP3ZufiollwB44HJQKWAtOY9wLYW9ZgmZq
ZWn+l4pIsJWe+w6VcuFv0uPljS6LPaUP5q9aCTxH9JUPN95RC23bmLXkgwtQfqi/82LdQj71H7EU
c0CEcUwxo7vPRyjUQYN+frp7NGUJyuFeHU50R0N3PLOIzAiEbmQ4Qe3X93GSSXZBTzl0LR/5WxlY
iWQ+H346U35R/GSRA1A8F8QsTsV8upgReuosAnFqFswfRLn+pJMc6qBwy6F+GWpuO5BmmELirz6g
wh9iaaZ7FroQ11PLW3ylAeEth+lhz3dO946N+OMCqupsWpTXQizrsmRXYlNEaUPu0raTodHzKlOI
8yFyHmCz8ZQycD2nESusJRwYSI8OoHMmfVcxgNI29h8iTsL8JKNilXPIDyCtiFPGkqpOeN0q7JXq
tWZigIvRX/97lHJLUjrM3pAjJnYDlnovY8/0z+/Nbuy6Y1HHkEAWQ95OnxLrdtRSj4OcVupgnV9T
7qk3yUKb0KyNFJ8H26I66zd9WYq+q7j5FoxKEEx5KXrnQC7cPxWcV0rQcnRJ/XZbD2+jLNbqAT14
K86igr9xURhhrDqI73BfYooxs7FmA4lvhb19GaOM6x5WkKXyRbtOesv6QTu33UUFbg769zUfCsRy
ooAZw477spCuxhU/hA1IwtwUq95/XI1nE1xLYHeNlLYZBP6N5mMNcA0i+h6z1/8xv6BVlkgt2Weq
isG42nwxStT5VfaC/n2r/wNhtgPaxCV/3O/Q3NSN7L6vzN6zbPjlmNDGpUEWAP7v4EVdDX5HPxJa
EDsJlIdRE/R0M1omd73weXbIPWTH2Bfudz/sabL0iqcmx65mGKHAAlDizli01EF133+TQPZtiuTl
+dizcWK93HROTPXh297WoJMzmpaq1o3jry25cyY6yL3oEWzzyF1TK2r0ngfYNP+LZ3fHL+6bibaK
ZbtZYAtf/1CtM4ww/pfFlPuJ300uS7vURCVmNMY+7198xycxrQN//KfWCBHV6FxNgtO/eiKXxiKE
bedYt1iM+NYOw6p8KWMUvD63WqfUUuqJtbC2eYefbmQMUHf33h1QlGjuZhWpcT5jsI18zIWSsZ5x
7MzpHhuo/NrR+U3ZFzuP70BqZwFxaV8CcXhQnRSwEJOKXEc6G1YNY7WQPxdwtFuKGH8dstp1uoBQ
7b0d9PbGU+lsCFhCzjLDvq6jN9zo3BcX1SIXL4xtr3bZ5Wldx3H+xGtcKjlbP96H7AgRzDRDz1Ep
VbJ0l1WsttL4Z0SsL9ezVByEhFbz2wqRqR6jwNFJImHxOZ/sJO55J7QQqK8W6X6+Vti9SY4XuPdv
kya6mSZnkMv5V/Zwo8QaKxEmD9rYvgOIeOpdlU1PbCueByHA0P234fgf/YOlEcn43axe5O+XRm9u
GJm1NRjVqL3vAnpcH9VT4OTupnAXh7i7ZenWrzz9YzNQojVWLa3GWZ3uRavPPTEpCmfRs0uKru2o
ju12Robgc0GSOWtVnTVmRJFiWdcIpWABMk+PecbCB+IvNuGXjXnIiX7NA+AQYwRFiUrC2KxfnM5b
/kG/LRMuxaz5ZoYgLXFk112E+oMn4PAS70Ah60j7pKAtrPs8TY+mInlGcwH8XhBzn5TzpPiNxJ/e
31rXmoj3ffwyJdJO+i76HrTXcHZgzx9SVsg8woAWMYrjWDzoaii6v0gjz7EucC5NGYsbXwQMeQrk
GxZKFNpZZal/rK7CXh8RtzgxQDt5PTOegrBWDZ6dM6pI7Luuz+rIl2/oFREJRcMFcgasR8Hv1cGm
D3K0QLl6Q6cIKVRXA0UK49/e+24rZQLXQu7/ZUzN9Cr7ZieIlK4A5bzT84GRt5hOY6oyTIzUiwsg
Hv56R71sr/XMe7sUl79B+Y0QOeOlGNbsU0lhQC7FolZOmbqwljgS7ftCo8o5sVMLh4FR/7ZZmG6h
uqqqYJEWIUqaiDZ9QYff6vgUb9Vixryi3ZKFY81/2tZpFihwOO4YHuBeuluGpHr/CNl7TWwsEMr/
vsWuTScBqKKcDD7YPQ3E3hNhpY9B939o87sFhtlu8tEbFh6i7Qo2iWkvOYxWYZ3troledJCNN5Y6
4cxrPigWkZt3DfkZLMDpM+zuLMDnjDX1ujMywXmE44gRPSm4LTEEeHT87b8TQSublrfWZhFfNZOr
7oEmbH3iBXOmAx0HnmCOqzlUie/BiItR27QHbT1jPu39D7XmXFFAiQTtwsDznyiAFoxlsFXobKiz
4aAXDtGWK320qSu7H/d0mi2RIC/s3ODZhoy8SKCVJ2kXH9m635cAIPNnXWUFOFfwhk6+s/VlwV+X
52vQ/jVoCpZnJkWYiz0HLwj+ku7pTvbQYIE4WmgPkA5TwS15NpeTSueVE5qTw10HVl8R0BN8ZpRv
nLZCiJVB/1eS6VyEJCANRAdK+MAlgQmnUXtYfvg/aapgcsc03AGpCTKS7hQllUY/gbaFW3fWx8x3
VmKtHa3ZfcAZcNIH0zDT+J2PkOLfijislAxI00xX3f1JtiFfNgsuIfyq6qfqkvvXLuyzISLOMcFv
1kXZfIutpmX0FR+2Di7MKm1eHMrimWnVwbw7tJi+BW3lIuIhuHOAU3z8+UoJCXtlV2wLJXR7INP5
ssO0Y6hqXfLNc17YV72WdzGFLI+8CP68yvaBdKPdnwyhGzZRUf2jRuAaHJVwelwuVe3AA/vwyUSl
6iGzZX9/fN0dJ5BhaE1z9ycnN8hok/inlPXcdMGQKpPk+sLHf7VGx+STBhYLUE2pLqPFZAMy6gFj
s2xO/d7OySi4FknU8uJqEyW2ygIpnPyZjMNDhXgAnUC+VeC65VK08HKdCa6xPC8gAKmcQuFuPLdd
Dzew9hQzfvDp9VZ3wpXf5k3f7ARDWlxn27/0YwSZ2pfWJB5EyFJNzv2PvjKSZsAmLf9OwrftloWk
K8Sgj2NvBqpdPmRpAzNqHcB/VuSu9ANvD5SrWCevSQSHjdfTcfYxmUQnx1EleLiOTOyxwBPn1d7M
UsKq4eYDfszP9xknGKxFpFh2PDB54aXm+4G0K8n7uBJN2acTbeHjSlk2LEYLmvlPTCwfNKO/z3/P
JQsP/q2ieE4h5NG6+ojOrFxzbP2av5BUwMc6ocsKDh0qANw2jSkMj9pgmpCe86fzEDWOajiyxEJK
kk5cFVoywXhkXu5Q7I2gj/kdXr5vLY1WdMPKgXMWLWo7jr/XKez4pwAy8zp+90cb7X2jwsksqjsQ
9j4fAF9x4NQOeHOjMOOcEYPg31BuP+hI66ZYULqPOFR7+x0/nC59kjACE1hBXsnaoAP1xkQtPhO2
YMk7agOoiJPhytKNjfmmiL++3EYWHBx4zaXCaEtt66fvE521CPrBILCrMATETBTDCt+xLe2dZsPt
JQy73VFI92tovh+GqiBLocdnNIydE8OBhT++XteFHyAej1ZQ33i4PuGa7PcRuUTaUd6vjaaaIlx7
VAifswy1zxhbzaKa0GorUS4l8/LxF7+R/apPyXwZDEfIzbqc24BuKaeDGRxUpjWQ+7JAqaMJjCCD
KPp5yuuHyCnRwi8qTesPMVDn4P8FDwAprOmLuo/93EvGeKGZeg1PDWnI2rhr9sgFTRAnI3SoA0XM
3Eo76TD+82N7LgTgU8I79AM9BiEzlXT0D4LAg6VI5C6JAbYCxKpLvbM3oJqzkdM5mpRO5h6McGEG
ToBocAMTX8+lfec3M5od39BAOoqghdFuNNN3piU9bgAEJcP21RciZ/wMxbhn16JB4t2la+ml3HGX
R4loyfLyON5HTyCYDgxO/1yb1HkzqnKRCHpVx7oaRx7IE+kTLodW20qnHkbhQl7yv41AyhvK+jIJ
AiWDaXVuwIytjeFrGu7AhXxAN56JSplQ6TSwScLG6UtZA6+wvPqbOJIx2zcNfVaJ3jTaW1eCfjOk
s/ZdkBYZl9XVQtG5PjwfIyVi7wvE1vSmehfpAFp20AUYXmP5ARUa6y7oqGsyp52N3V6mZw+/Tb2O
X00JiS2f6yXQDJUHqhKj5wdiAb4oWmReXl9mE1AhnrfjVlsQHjZB9BgMBhNRqffo67MBzK3TsZgT
B3VUHaqaZaIc6uY1rhV070kerX4iVTiQZy3i6BXtNyNc+fjli/BUT9jTFD3YjxMQdn+xpd+OKZDB
Z13dyPdaFWupyODmaj4SqohXmjQuHCxQ/cvyXacV6tJv2iY+D8oNpD+S20bGatloxG9PnI93SEsz
b4pr3+dcY54k0iNP7CFRsRv0zWM8CziXteaY9DMrA+UncCTNumVJP0SsTqszOog7P70YCDBIv4cQ
RcmiKvtifvl+kbKEKj9442iuBCsA41o39aP2luXVzyPoKPq6I4gWO9Ds8hlmZfxV7C8VAiIXM1EL
DSJtW/FH4Tb0O36+1xFC7qt6CY6/0LoeaUH7KMIxMIpzvmoI2epSwmK3FGbBqOUO6TQXVz3z024P
EZWnXNFr6LL3Rqdlyox+7+D0OeVvoym3F51wDBYO5YYynEYZP0veoKVF1OWtbMsteN6CJ21KxWpX
QFHc5gDgXOCq47YnddA9Tllx68tYpAlGimcHUgORnYnpQNZhVBjwTraAM6iVVH55MAwhdKFdTUdz
AJRM8qPp21ZqhsQOGQ9WxZCdGaxpLOcVsHr+gfE2kBUhtyfgwdGKd+RVfJ2Xc7FA9IFo8qIeYRg9
FelPKkYk66aUSFx2Z1Y6SCfj/bFinR3IJHk97ZJzsMNTqKYv0Vdj6pf+EboZpBPVE4iPyrd/x1WM
VW1l2J8EQFS6OyUDbEyEjqdKeVieRfTrys4i9mzTtrjCPP1Tg7iPHnqe/VYOrKry1lJvkJ3AHm0y
FbqzyMA/3fQNOZ+A2oc1ei+ezHyNg3s1BhqeoJ+WR6y48dNwe+l2DNwa8LGaWeGcdEGWHHLySaO9
54wDnUCWdSSvTShmkFDfD4UsHQP6P6ZGpGF8H8mgaUsMmNRUwAl4wkhofBpMfVVEyk+qbQNRqE0h
wMgfJ5myhWynBYxsHSGfRcG/HTEnr3paylOHxjjsdj50QZYkiqJj8ZQ09r92KaahhIhKchu2karn
murlCcqA+vyk3sWUTXi/LthKQjnhNIrOrGF3v+CvirghWEEBgIuQEZ8ZEaTkMODCG27/wMROJtoJ
R9v250nJ4e0yc1Lv1HHBRda9t3+xGtq7VR/XkZRsvdwOyhKX0hX0HZRnifuUrf0SkhHrw/K9By8o
qva68BOFrCeL6fWpRTqID9JZ1PQ+6hx/TqueaNbgRsOOEJ/hnElQNDllJzM4HgtwB4tHd9HAbsiH
atr7OLqylnWu9qMJ3ikSkRslJIRnRFqldwfSnR3+cdgwFUc8vaM+C2+yyetLDEH9qYzqXuMLtnhr
bY3qWLxbe4vWVGE16V+cV2BmlNu2aC8JVHphC5xiOl2RAnt5qBOaMrlYHGaHEh4ZL3+/EVnCxVIc
8PD5FZrDFcIOfOKLCNwrFPudoalYvoBGwXJQwyWQB6xxLieyR45RAQLXuerGxpSqU1W5W505n4Yp
XXAkjxpYMAcV/l1wrSuznnZ1RVEiyLGrGy/Fr4jKELSmV3+L+NMHv7psX62nC67PL2ZC/M2MqFDA
79rBkUpC6GAanSC4Imj2FXLEFjoXMrznaUkPgSnj4MmK7MPnS2ddMx+2biazwz2z+buFt8ukTD+Z
KrRjBIuhyr1IOaXRXzTkuLW36GKKzRdtKN/+1N12VICKtcwfpPSuyvGfNITFGri2PzIO6mFz80cx
X0J4H2T5X4WBqtiF5XM3HqqVqhy3sxc5kyI9EmzeaTWeK2iDw6ktlBwbuObuJqax6zw8Uy20DSwJ
ND7dVXl0384UX3mhjjlqWsltWFFmNss+9uR7A5r6YV2KXInmULLSUZoAa8xbkEhcnt/u5DmeGMSC
uk7OtVXNagf4QJJtg3OSCObSk88I6/H7gyvMQ7VL8wDeEW2iIhjQa9ZPnL49INr2c4feyO56+jvd
S6vTkwRNwvChaGVD3Ju5jJjpeg9TO3PLY9IQsQDAuXIo80VRv6BN2/t8NWsdnOE2bUa6YqQsBpE1
rOICKPFSYexWUCN9pa5s2cABStLKIPtrcKk9Bf4pNiTENhaOjCHREA/JqMKbzldR6QRrw5tHYbue
MbgL8qPaP49oOOUP4g3PxEZ41BOyzzKYmmt1NQyp8Ou09FLSg+RgZ4aTcDYlxyX0pqSRGaTqC8ah
eeoy7W7y+hWr8/Gwa7zzlyK0HHX0HgLOmxolhW4P6W6wubflOGV7Q50MULTuwFeqZdYxzemPely4
hfWzlOhrWGSm83XHcs2xIsZHvjSV84vocyr/78YAMdEnJU3yvdDuwe35Ci2cj7CgEraJcfwtOkXl
WaAOIIAJ3egTzEXFzLty/eZbnmfGknahvC0fSSTGU0q1sfWROQR7jqmG7vQc1S91AZjrW/YaIiOr
FTPyOxzXc1hKyzzME9mI2gBFAQfvNm5suDnachbRrVWXj/jwVPZPiIvYeSvgTEjSYUZf2nN3LswE
OaGxlL9yFg4FaTtykVJPN3UJ374MZL5QPPwi8t63V/dHX7746pHuOs6yoPt8zlB+Qjunn2IIzbeA
wICdd89idN1cB3ousBdQu6qhyZ7MLEechF/WkmuVWvAwf4xtgSMYXFF36LwbqAbKRdqfBnD8XL/O
tIMJo3t8uDpEzAM+cGpaB/Y/46/Fw9RueJGn/Nf6t1kLJExMqhp04nKFmwg/E6YQIu/+UWLqHqwx
ls+CDKc15GuKYHNtFTvpT6AlrMEnxK07I3rHL6F9/+TTZtTMU6UIqA9ulDnPBDFG/THwCNB2z2Zu
nS90YqYnBCNo0O0mOxUXACOnxQL67eum327Od+3Cz8LCucE9xQ/CWwE6z43/8MvlAXXey5BtVotJ
iTrMtcswo+osXcMUZSghZ5RdnlkheQ1o5PgAVy+nb0Ofpua4rZz4S/IYcHs81W8yr1K6xzXCUNbw
bsAAMwnjdRbYnQL8pus6kdt41ZADghaygN/na66XMzsmL28fqYzQpsRDMBTav+jF0am0Ksm5ykFS
fFMBAPOSEaTXwNqanNbg1TobMZc+yIyU4VtMXuWc1XgeciKmy8xyHdZU5XuvBcmBBb1fA68mG95x
eoy1ynFJcrSKEcWsgu1lkAw990isRgO27L4/TB3haQib5PyFjzDJKvF3AXpE6kjdFux8KRXYnvtq
EyuWbV4VVczXXY3eq2BWByx64fGoRL7WciXhUaB4PKH8vPHzDPmqsoG7DwJr/sT2Hg5h6nyguD3L
zMlarLQ6azysphEC/e45yARX5pZjwVN5BnswZfTDRASYeZ/8I7WkcVqRDjs/SpZ+TyNofN98XmAz
WDkgWilu/cZc0ilrSbSBkqW23vUt7949yAyqLSK+zEeXMsHhzRHjoGuF0bF18nCK+Wgcr17OmqQt
rztn/G5Xa25mYHj4hbFXoeQBptplXoz/HpVV/wg4R5ZRuzIJXh5FNDHQUH6VWwIh0rj4e+kGKaL5
4cXoexRG9RwJsNQY5+nAytihKwhTbp4OiBQOVJPbBCdbgeoHpLLzYyNDLFRQXLzpMgCpuTAL94LT
TfwxbzYBWqbV9ixWWjqjPAnWfDAIxB3SxhzUuz0qOGOfKymunsjxlXmTyR+hjsIno7/WhK3KC2pE
h+ZXrtUewdn3rQ2vYJphiHA27E2ab+5RlBSzQGUWgz+GVJOXuzGOds+08J2cBAc8kZhgta1xSOVG
vcffpWMnXRvppO5exlJFzJf1ZAw4tkZISZxShA7i1pYn9RZdqv8lTyK5B4WlU7FCeDJHqikwhyYU
coRI8N/+jI2T0IKKUCE9drdWVaovX+1UYzsYs8rldmLzewwVxjPzxQjKuw9MS/rXqR5ZPtdCkxrP
nvxFKSLwu5pNxaIF/ZIMfTgfmNjRy7p0lCaRCUo4W+QfDsNodZUgm0ErKMuxhfe3AOKMionY/UmX
T67vQ74HYIp6MMiV2SohzUAgSFTAAL9vfozUVTqE3AQ2906Zs4yc2NurlCETq5KaQV3DiK5juxE7
CEEnUw7mAexhZFwaLL0uuXxqekz6R/zxvk3TkPmCIWLI+DcwlrjtuOC3lQjHYruqCrnX63jMZdeF
4dEowOXBu/3W8E/1/YLsqnwmG6acgQEL3V3h64VGz/3MxcOfT1bVlPcFSxbiVazDe5ors/vDPqgf
WVfpKtNuBs6ha7mC7xbc/IV7rFAJr2HvMTyttfZAuzSDEUlPcH5ru0d93AftX5bomAQaeUdYdT85
9/R/MUlrnNI/HTRi2+mxrKQQus1dpiHWFgHIboORgjVo+wgbpzbe/HvexqgfJRDnp9tT3ogZAzlr
Yywv4QdB8a0ix78G1mC7dwNfC0wECxC5YHQBEijQ8wmOrNQqo485BDVTYWcyGaCZ8hC2j6shkbAX
BTi1tTvXQefvpTNb/5ymHycGXJ8Tm2BlGly3S+BriyVNCdohnBB764Fzesn0mQKFpp6Sx6RhKw+n
XrpyEBYz0jLW1CCeCI22vP4HQu/UxEiIxluoY6v9KtcSQOlHEkPlyR0jyARqoM2yv5J2vdNfeZ2a
zRxN+XacH7QZlbq/gDWtQlVJ/xFonR9YBTrU1iBrl3M/5XIGSlyLrdXr6u2u6tFSdMa+QAtqlgQY
ygUT9/Co+dZCI0K6WBVqkfD5+HDZH0nPGk7MibN2/rob1qUNsM154uP2Vig2u0qMGMQkZWZ/G/CZ
mqjO4/pbM5OHUhK2Nz/+HATvxwkEYMMvr1NoG/4Vyhb12eQCr+RzgqffnP4zUxWUas3mHYYbJzJA
5Ze7Qo19pR5Dnc7xtPJa1Uq2fOsj95xA6Eg+vRCzqq5rZs6AlLDTu31oz2Q9umVCk+XR4gKOKVP+
2klTR/0IkCEMEtaBLd+JJ6NCd6EcoO5RkHzpPZWR5rsjZzTHXGqHVqToXyG8vDkzwIay36zWI8FV
TWQ8qxAecHLaUExbSypbtLcn8FL4ie4rQy6vkIO1p8SqefSawkDcgnmiiwOikXEFtdMUM/FqzzeM
06+0GO2u54Q+i9eqcAvv9ABfteIfWyETKGWq+Xtjfe0ltd1+9PdaRYNMgM232VkiRWJHoor5qcUs
ZK4Jf2+skgbXvdVOZTUv9Ag2TuHHfaaIKLUNXyKRFMe788ejcq+iYYhfAOflLPCr95vtd5haHo8O
dRpf6wUL/9oTmvqVjE4sVuEuRbM6O5zHMjwjwEznwlYFzVcupI9+LUNBP+rVbiJSQig3jHIQjkhO
Cd78GJ020gCPZZQ9w2GxYJ1NNtQwTUaYymK/F11HxEo4qmqaXNopvIgDSoAqceDjUQWwL1V7HaDn
h4VdgkH31EI35n5SUfGf+d7Cz2vHBrL4BIkoo4Tpr1+GKoanlLV8OIVDgSXzOEA3hSlx8SVQch7I
gfogyAQfvwSQzdP8CMekglZUKsgJiLu7WZonvHOEe0MMwhuYS2E7uIFdUaYeJd/k3IuncDYZEtYh
wjlKBge+K6jgakdYyCAo9Ea15HdE9aSHw6gPPKLWznhzfY1exnf7d662th2IYy2l/1P4msVsEsrf
3QFynx9b0V6HRjfYhLeJ/IOkNY5fEWZsHSRXVKnZRVkqFQORwsmi98DeTZvSTKbcN/YiqYNcuf2o
lCd86PjPX25dUK/OlQEJydsJ6vHkVwdgXY9Vs15RQHMI+0++pEvFy1Z8KbMIB/rahVJssPntUunR
RNFCrziHwBzrYCDJQnW3aHlquj/cqljcWCPh1JbU1zvXI4EySwxq1sPbSVA2glDdoOPb/wP2ALP3
NNYIP/ilCEl5jVneZffRDJjYLTwV5xjA3iXy3u8bSxDjo9j3R9vTBEMGT2y84yU1oWC3IISJazYG
LEX0WvLwJs8HZfrCwjGIjhy8aowx8weEwXkaM/0xHROev/EaFHG5ptl701oMgorCSuqYW+A9Bfp3
HcOGmLLW5JUHGil1n+muFuyw/EaF5brpsWxD7cZ1AVuDrjMwtd6aseLkbisG4x0g1XkoIK/xJE75
D7fQX6L+EoWaOHG5cIRiGKu6M+PCjhUDfSulWtv1FpwAO9iSL5/LDcvpa9aOZpcBMoYSy2tTeDJ9
KaSXDsOyapVEADXbtjkzGlkuJcC2VwlL93iw9bOt9uDQOqWtrbzsEUW0UkfJk31RdDwV3RhxzmLG
+iuDTNJHqPcgGqnHuqqzhbFIr2I+3SOOp5cxBOLCrPVgjMqm+RbMdsvpRd1+zrQyDsqbyOGuzp5R
Y/KvpUdbEs+Ti//7+GzUPuWDrME2jbCwT3v9g9Yk2wFg2Y0KnHHIfnJz0KxnfhMHPSjiYSreFuCV
80ExUCLUKBSdMMJvHPaxZ5mbkvisqv5m+WietMO3fuGjvlJfRK0vCivlUUhcOQ2y7nmOn/MRrsdS
YvkUURGay7iHnvKLjr0ZTbXt3Y563W2SlH53z1BKq/uAX3MfPHVSRPuyCTlRYSYUFrkBOwNJzGh+
LlskdGYXiYsjEQ9ozveoFeI+XIfJCl7HnUjFncpVcQ3FGbtbtfd9uxNYKEYxgzXvWlWnsEX2H2Yg
Xy9VnLj+pqLP1mFY7LyZjVXycg7RFZGFft9x06CozhiEdz0OBhfJmcev3vHQs5QhHiLUPOeV17ow
+WrPkxfvCes9zYkGlfsTo9mppYoYH4chveulZcKnPw6qInUDqG0P1r0CRFw2RfXsVKAQPRpCeXcD
DSD20t5/W24JcfDHKvFffAoSyetu/pa6OA00tdzkjgGCxwyTE4PWqvTYIkEvIqnbMiBN95aN3kAh
TspVOwuFvIoxnodFWyDJf1ySV6lo/sj6jc+9HXtsSIBglhh7yyWXBeFo69/jGGJ0f9oR0KZi3RPP
mzCr83vBWzetCgacPBMZp4hTK5UduJ7A5v2a3ZD18u5sa7sUi0Fviuj+c1ELsLFjS+4WiSk+1Blz
qNsYmxVHsHUF5QFG8CypHNwrgF+cEKkWmVoikHFr2Lrkt0rg1tk7QJj5Iq5Y8l9bpe4iA5rO62vX
+X+gSdao5bZyrBm9tC0T+yt9MTGU8OSTaj5x97vLd15wzHPPpWeqCzx5JUdR6hosxCQZCc0X0ZBP
BuNgjuoUYVgH9+dvP7SC7BmAoP5urCb2qnhU7B+IKq09FGkmcAJ/fB0xjTyIcg3tDOddonwjJclJ
i/OzwfJ2+k1G+lJZMXkIN2RqePY/NQfaqzoTcDLr/gvZrwKsgjmlTT2gqXDysLWLYXl958/myGq0
aztGEuQC+SC2y4BfSVTvq7CpAnJ83mIu8sj/9E8r8pJR4UZ4pgXMiRSZqt+/dO+ifPIAjBSGVfjE
IrLffQGBH3vjuKejJdMWze/8vsGL/Q0g/u6BQmRrmJzxD2Mu7gnFPG2XqftNiDu1+slwTCTPTMrO
GOfJ5kltUp5MSeGMLkMJsBshQJVhnaY6K0AZnt0NZ3iytxZkKOrCU6o1G1EJ7Fmuh+Zrr/FTALUG
L21CZCnReu0uiX+cY+K1p27Uwdfz/jYff0a1lpURRF79/K/SybQBif0L5wyH8lPnILvqxyZuQAvB
iP46SfcpdFiKO9o170SWmrF0a4hQrbGYVvpz8SJvW6Lhfh2EvwgmcMoadafmtun31gI3bMDqTaXl
AZXuEoFayyUEf0Bb1Kas3dFKlshO6cvtVy/i3NiRRBQYh2/CjfaP7XlW0a2VR4Xorl3ali8Xa6x1
VJSpEiKFmGci8m5+X7Ig2Mc9POomYAY67VrLpto8Te2WuKZtAuavGHsu6/y1S4g8GQ+tOGfN/j8B
87489NwQbbfEGVSSCWzax5aO63RujixgDFB7kJ2/aVKwsembs20yxUsKGJcVf5IDuWlkwjcTKOfh
S9DhCyCseRPbbyQPwan2on9lorHF7B4F5wbLZ6TTBRFFK7pWeBdakN7lURYK9S0BjZr5HZ4pXfff
AA/ZTTau0gesdp3DsZ9KbyLpyQBb6ZEN47GHeNix+yhYx0lDBmf6m7MxuV34tCGBtx2AvAXxD6yS
YQCSw5uWlqhw2Tz7t1HqaMU6ieMxCT9cvE+XjSn5Fr0VGVrv6n5ubsfj7leLjJ+6UGJkukh4rdSk
0U9j2WMGGU0E8ZorNPlNG99xAyou+F7GbYa1QfsziuHxiSEUluYshe2IMAZ7Revtgj0Zm2pFCC8V
//EllnmccOltsqhKyvz/WNgmWeLhjcYHPxElBdhzV4/28XQOzTIMZO7gXliZw7Xbynjn3NrQZsDz
QTHYSGQoNnv/+TElRMUzf9/l3+tVySKS4n1hxbJA4U70LI/BzTus88wUYT5HfHRvYbeOe/LOgUIn
2fUkAGM3aypkRvDO9aPtcu4OCUdIEpoerQKIAH1uHYHdx4KL90K2MERRXXFasv/irNtvEkKmJE1G
vsJB1pqovmpSJ+VzyxEkOOfZTvY3do1VY7GIl0tMgxZKNdCGd/6DvUdpsbuEbK1WuSqN5PhKL5lm
pO3pgjgmiw9DcygBHFGO8zwdj76b6HL78wHt8BANk8i2YrunLY2q8GvZ34Yj0l3qHepwPDYTZFxy
IygADNTIlwYatCJlJ/jKZABanu6NFV7b8tMUN1xD8pqcx14XboduFLWAy3RHtm6lSrSPaLCOPstB
mOk+EZPP7BckI3Ho4Y5SnydsVq7eMvlnDxnkq4wGSR0qUqXKrXYG5UTVHJiFOPHFjQVFZlp5ULyA
X2HBFnUl8e9TG3dBwK57SxSsgceHfg0El/Du0xRWDEr9GfEE3V3ECIVrqG0Am+R9BYT08/dU39Xe
/L5UoANRAVoEHLLvsJNT++Kz9WlhGFg/exl5yVFGPPyUgD1JquspJZCJ1jLztitQpKP1lMCCV2Yh
NTDQUveeM4XjEw2MR0Air6mUc4Qz8uzuPU55iuMk+p7yMEVraaCkSgeoIcdM6q12zMZxidge398T
nBL3EZcp9D3+1ao6gJoNjr0En8QCSxJTWABwtmOMHLG2BCgj3Isdk4mcch9xDOZH932u2DC0P5+e
FdnjBlWlRx4CfdH3Gpg3ZHs93K7b8HhK0YtPi0QnIPaulAIXhGe9qjgVCYFjmZKMrS/rzlvxybLG
rln+oMBUBafgloeZH1SI+IjEQ/os+m2wiqVhT0gX06VdQgRr9ad9+1crITJnrYd9p0o0DV94ufQ5
i4/IxgJVEg1jJJvE+h+w+QLb7CO7njwAO5QwnsFPffn22PAmnQuEZjmffm1DFUcvgsaYIokaGz6E
iYUqIcKRi66hmD1uNEFXkSji58DtIKizB6tGKvBCIcFFkMChDdQPTo+8rl48oZekrfuBG7CkVmv0
OKThcHYnw2EUxhjdbDDGXbjK/Eht3HvxXQzS2SwLKk5ofqaIhyEPuF4LlU1RZGuXWYZ7eZkeT6zF
2XcaOK5ndrrM8A6wgpdOlSey7meU2et44VZEoTiyKrmt0olx3q0ouAJmYeBV4z8qe91CR68Dvt5k
xhlhjcchfAYO4cvmIpq4wrIHf3CiVBZbeSjoJxI61rsg4vkoAhH4W3BQjOCvG6e/4u/w7WTMpoOP
nu7z4lYV3r2KMf2fdYB0k6/6oa+6M/ozJHYtx+bqlPZGu8N0saYkoeX+rrktHKiafGwjFHrsPc6L
fZfgQ04UeFVk9vOblcxtHzuUK+a5Yo0Cbaa4bLZVjZ+OdwLMiBbTiYoUR7a+6MTwtQ+Dfkhh/9Wb
gKzHN88nSYU57ToTLEfDstbgeemrWbQ+VBq+dxfYUa5+SJW2b7YCZVQygq+XGDLBi7wy/dNc3dak
Ttj2317tYgy8mDQPcLl0rY/q6WXhYIExc8iYA46z0W8sAOVJVXbwsHwWTL4b7Dy3A0BSXvEw5tWC
TopFnCGVaWzVdGMjibsHrnNUsiqf5Pk0U3QXt7/2y4NX8Ntg6txJoW45nE5dDKaTuj1i47SDZCCL
IIepUGkxLj9K0JQiwz+57L5FoePSGcV1jEeoRLoWC0LXGIbXj5CfEC0dot/p+nS2bgzy23eDyIC8
lmd76zBJQjUdTCyomR/5OVKujBPWX0YdNZJuyqNV7QmFmDARETJ6yb5NXGlOHiWP7B4w3tScZwWt
xoGl020w4Hi5fSTZk2g/UvowjZxWKRhfcDvFr4+6ypyedbHU8/shye/kD+oICKQZOJPAkB7GkSKD
lDxnPrx8NnhwsBd8hpoNehqVemWxdNFZHzrPFG1C43Fqn6zYQGUqYVzSgjuxHqW4tLHYA3r8eTTP
TQvOqkZHh8lKOroYFt4h52eCTPoyBznqTRU7IrTsZZnF+QZSY9JeehM3fuXFeBIumlL+67C7Jctf
0r7t7SkjTkNfKY98FtzBB/MZN1VVs060/EfsevX0j8iuXTeKJBOcwKGnafMWIXL3C5Sg6bZXPs7I
uhr0FmqiQF9EK1aY+H2u8mOc6q9tFYLI3BOmQB3Txkt477L2UYaGFNvGXnG40Boygs9MoYF9v1f/
2NT7AO7vT9qAXHcpx1k/jQB77VhfYNvXucwUQjeTUk7/JhSgRrqztQ1NHk23tiXUS151EIPo6Too
93o94ZzXIj2ptbcnwLufcg2OD0VPBqtcjDmf0b3ZW0Eld8IhW40f10P/T3EnWUZBF+s4wp9K+wSz
SDfVWvq6Ngdnwt0FptKfzaWdZHrT75Vy7seBUjtNkiK9zGeXZjLUG2FbdN2JAOwtlOr1+q3yoE1/
hTatMdPh1VNgkgMsdQo7IJvVjI+jtF/oNZuCO8sORfc2V4Vyjpid6BZi/pjTuVSxNqGZ7R1/ZSnT
1h+tf8B5pyINLVfzp36FLMRNAWZAJJnk1U3p4J70UMwu7MLNOdsJz16koVcSdS8opwti1jQitimX
8rSmDO90mWE5/6ysaMleSH2aTfWtH4Lbh+du/JdqRLb4FtQbipa2OA59NdokKUTl+3jnXScSdw2U
5EUjg/6DywUsDGSoBIentUn8erFI4CHhOBaYuJ60CFrC/Jio7gU0Ls1g6JzGnsmlTDs/HUoP0mC7
4f5msBer3lHzV9YGO60f9yk5FvbVneDVEHzMHzvMPqvg8kmGvgeKFt0w6ovEuyYnMHFCXHni7NZe
ne9crkBILFDkkn4qK+5frQt6toU2A6Tkclr3iFYcuvSdVxK35m+TzgyPPrQkasHhSlKXv6y9myww
5gco/ViMyBvyjLTaMTyPQ9knKxcZAbElR2uMU8XuiGONQTkT+CLWXmgShIboq6kg8JAVqOCVHR4u
aj76lilhv/PEtrN+zdBKnVA7OEnMrUhEe0+yuEdCcMNf+qHlUyPZBa5KcTW88+eA+TzwPdqwrC3O
ylMqZI1hBOLtX8bnGwXlE6piHVjteT2+hhQjp7VOJlGD4aUI00FD2CNLNHl5lhWPeoCcie2DS/SH
BJXn9eRSo3SsrruD70ClXPdwW7qOfkpTnTwg2qcj/k4veGq8DyWUJ8gxB0Z8XbPeTedLu8kUqPeh
uWODZMHXNag52uiGS08Ue/TeJ1k54XrsAMbN3rBCe/rsRxwS+nDBEaosVe6AcyZ9P+A/gM9OBssd
U36w6kUZD2nm9fxQ6F1iFtOkMkEB7WeZxqVcDHSWxR38FP48aOmsWBo5Nvl9VqpR5YGITFGnghDR
+p3fhp6fgLT6m90sNAoymYDzJ5f/Vg2DsxoAO/JHgdkWXHEU2FGDF5j72RxYL3wSYdhEYgKkwyio
Zl3vunzYFQWAx+heC69QTM/wSm5SpNM5sifyfioWV6z8nZY5g4SyuY8hXdzHuFFLKVmjllkh/cKx
wYrT8nVBqtn+CJB6/EdjYTdILPywgMzYyXk7yGlIzvLAX77h7bHcuymlSfttTJCazO26HMcpfL77
HtJ6y/QSTP7tyoHNJjRKrgxRX+sBSvVaqejhhRoMbTVBvQ0zfRrt2H8yvrjIGZ5Am6V6+9xrd4o+
szs46SCZTSp43XQ5i4GHk3Hp8BiH12fYcBo6oc+imbshtLrm6hq3LbVyfX1QXekTJ41uas5V4AxH
hBwelQBCjB8YXEsh+kiAmuVuP47gkc1Oo+uQTdV58g0IMYZSO5KCFiExEF5XCMmC/wMB8F55vfT/
bDvets0CA11NGPwztqRIY1JwxKJjfNroAl8tluKg8iZEzngXo62+1B3j2q4R1YdDJ93FPwqsz0nd
3O4H9eRhJYsQ3Llr/TS4iR4+1KqzKdnpyNKq4omYE+H8cO7V8Imo5qBeJ8CUon/4gvpJwjj6prYE
xib/Hv+yiOf90cbM2u6oYcINDULBXLzgZbe/BXVbWen4WbS/TBa9EcyEhVDN6xlYsopiCknxArYn
S9Qg0OAoYnjBMwZSwZ6EuOSaeqdymI4K8nCFMDR8rHRsdLhXmIFPnRKmPqg0O/vQ99Oz3QoZy24Q
xJi7YAWbKAYeSTHjz5+OVvE//8vNdh7RZzWre2DKC+UOsVonl3yTp/jg3gJrAHHE+mHpabcxb5Nt
YCcDl/abi8gYsJryiMaW5oXEQNFz6+pLOwu444mbv8Mg4l54KHhNopB8XCvE9xVzEEshn9xqbdUt
/8vD4ovadbCV/e0zPJvGKl/faYZ59Mz9NFzRjuC+PMcCL70b0u33vV92auI+g7fiUiKwNxVxMWsj
5bAPISrBxVN8R8myEehSVulwwrfVhfViwxJUFg2Kriham/8JSzhUuGVWr5QLVgKRT+HiODk/fCEK
EByQU/v9jMR8iDMxq+ps3iA3DJ/tpL6x0lyqjmWvAaGB60UW5uLjoaoBqQWx6O6HKE2gaGxLu+R7
PjswDFR6J1/chEcUFaM90sINYZglMZeFPeCXOIgjWPxj5sTakxzi156iHVr57fpxCHX8C4KLsoaV
pGepFZWmBr2bMagd3Mk/6ljNFP7SbY0v83lCcq2qcPrCfmudq0FPEM2NhRjIA/tjFG4+usIAbGK7
+I+cKI3EROGg1GEvnY7LPWQQABaGsdkonxk5EDC80JYX51NEVZylEHDIVntSi+sf1xHT7Tzswxbz
3fIlbdgVHLs4f9695/UpKl2lO+f8XjSyWihIQ/rKpRPuwKiGOBWNqDjtPOn3ZvqrzT8345aapBB3
7N04N8jfx5GsNQcu+J16Nr1+JYYgnN/eFicg+6FZFY16H4nZOqszpe+qYHc88WD6N4qSyNaAzeHf
gg9oEB2K8181svkg7neSqCDf6iaEWU0beJKKYVFIxU7YpPUxni8o/yOHx9yOQFPMk6ZHbuRnrrQB
1+0OuM0UO1P8vr28qOjmVKZhGaPbj5oPS1NxS34gUOY7a2TqddvZon+2krki/xVal3Jg3OgL3uAS
VZzM+RVIYLFOVgwAN5IKJijjFgM6Xpkbidv4z5uHWSR1vDhqriQf3H/wFJsCm3Kp6xWSDt/Aw7/h
WQWs1JirJj18/NzbGF/isXiUd9QvYzlWz31SROy56UXEDuO/tU7MxDrN8yksx1yqvUvE4yCuC7Kl
LOx9uZBmgT+yy9/S9rGuv7njpJPNQhO0OmCEYTYFfE72XodUMVfhPmi05f11FZgLKE83upmFNGgb
5lvWtbdEVwkRy02EFVTeWuk9JDoUAeDSfQTlNiLx/0/1DEAGQYLbFgQstTKltv03tRDaA5mQSP9g
1g0FXweoGTgxntChnpgj2JerGW3yuFei05rzhitO2H2K6HMjCGhHZL88xQ0oUclvzXDkIbTeP7KI
tvG+XtoGoBmYNarlcEUydAy7eufVm6ilByUIxNo6dHQPT35hjLBQvouloryoZxJCDP5JLnVJnD6t
IAE7mvUCB9q9b4OfOVqQLnBsydKpmz677mVg3ClKHPvnKQMcxS4hzuBHviZ7BnrWNOx9omSkAFlu
MCwKsPlt8SMcT1LV/j45I1WDt4+lUNnEScFmeUlr6xRUA2sUSaCdFF6FhR0iHyQwf9ZKBQNH4DFb
9ntnz+hbvYN7UY00YSg5dJKOb7nzqgFd4uQ17aCfuH+9b/7KYkhTV5MzmKCv5bwVjP13ojuBlYZ/
0mBCOaJxrTiHHJ7NSfr86PGQnl/ZZFnwrtHGfVmP8NLqBEvxNZVbzNkGced+MIlqc5x02W/JRJ/G
DCZ6W9nC4YBsugLKV2jfj+B7V2yboYwl1KhjaO7wpTN+CWPlVGCa1Ng+ewu1vkl4rQ20wU+7bvqE
RZhGkH72JC91zNIVIya9qmzq+QmKfUVZxnqSWbi9atksP+M5cHQaerg+vrn2sVOIJjo1NkK8TmAi
jcJt9WykwF0BgutNmnxGsx82iMLcKM1fi5UyPQ8+sUjbWvtX3a3OzxvcVsqg5x7tMgKHZoLayPfH
twJo9kSXw6TUM0hCEOApRzf/tS8fq1sHQ6CRUygHx3c9YXm2kamYSE45bcqXwEra0d3qajfoHOcK
/Yhy0xeBg1GRr8pI86EdPEZz/QgBPKPJFpsKIyKTjl61di/W4bPftPQSuZfI89q+9V2AKnF2wIX0
D5WhwaoiuBQTDxDhw4jd+LYdRzs6vy66ktCv71EIXMA5/Fjjk8ruyhrOjXo1sfRBIi87/2Allfnc
KNQGTUKWe3ebNGFxOTNOAi7+TU3qjBeNJFRwEX9eZPDGEDwOdnT736y8XC3TwfBA8XnWBJRNO4ti
QyyTaaziKLwc7NZxipupBznlyAQN+p+6zI/kEk/6PRKn2fiKa9rUN0REg/kdpC7K6deKuaalip+3
31nAn6PsK7dxftTHO2xpHeuFZ2GmVOsCeEuH4/+Ox+Lmklz6/EYZm7ZdORZ8eiDI0Umjz0Sp4944
k+wmgOKqJUhUZhVcK4yUbxPvV/zCr9GZT+9EuiOVnjw+rDcPfTig8QjW+aQLHv9tIQLuRH9moPXX
nsOkQPvITXIy0rq09OMjR7GItjJ7IA64sOklIbrBYn2dlUf06E5x1ss5Q79SMKkVmf8smiyYwJJC
hH2H+U07lulh44NusykkwiWU/COaM+W+Qgh500HKiHntF/7miybVuODdqeWYVY8uhi05kN4PHOeE
u/LkHz+OQyOurnKoJ8NkeIOLqQvE4H26iEmMbk8c0QjYyxBPFyY56Y407bACic9rsWS4/EB813W3
EWvGwgGSBNK3WxmZ+W8WNH1KlptB5FZtlmCrlcFMS1jjz5niDMwnSeyodb8QE716kaqAcz8UrL1V
LQw1yNdNGWTQJE3BGHQ7PLBPydAyQQ19K13M2PV2tIvQBQIjvOdt9Gb/mg1Drbcb07tR2i043FYa
xSYFXFeFhrAUpvkD9tpE9ayvcqx2hNeZrXDL5s0xUFTTEkSGERDRU2+V5qbjFkVsK13wmilfa31m
8pZ+4NFLjgR/VbG9/KX6Gu02lYNjzdM+2ueQQV/nNC7Si9rObXbiYqMkBOWaf1b38Yephuu1boPD
/DrN4+QQrSzbXlowS7awnkOTpMEvw7U7ULfIz69oKe8aJ1tom+3rSsFEL3o1gpvD3tw1Tfcu+qb1
MUjOjk6a13BDvyhqhb1vFp5DKnH8j5xc6ncHWlSD58hrIctlXaSgvmtJDST4uyw+2p8CKbuD2crJ
nfGIUfanwm2YTh2TeIkE5DrQdnLvm5Pg5ARrXsTSyrsoYFnaYg6pASA4X/MuhgsRiaDGgMhQEQOB
RwxyaUU1B7Dr0hjg2xst6CoHpaO8RZh49+sWQWWaqZqLu59FVcu4TOmAakpuEgTo1GN/blybLI90
RkuSTihGZX0i84KEi/Du+kNK9CzoZqGABD5as0oz2Hs3k6ALsNsjnqzRPCNvoBL/oBbX0SzqO3fr
7JEbF2ArabKrneemjL+3P3ryzimdeV0Hz1d4jIItImRsuj6IXH2Y5V4UqXkkB6DiEBZROAAcyDoL
gNTQkfuBjTS8WCeYhiE/o3k29Xp9xY7O+dbv4IF1UWeEJ+iNeoldfUEyeuINBv1hFfuGxK3lQKbb
SD9dV3asMdKmm+uIKMDj8sD0K7szk1hYbrBIiOOY8+Q6Vj6imqossmYvyukL8dx/DKxPb7ZgULEo
7fOgLHCQjL3AUi3h9NbLPXJ2nuL5SyHKEvU72TumP3gZc5x3Jepxct71Pu68DwO/AbWN9lplcVeA
Ifgrxdk0U0XjcgZf/PyMmNAXEOkoyBPquHa6nT/EozmdCoeSjv/nqCqjcBFqVD0XJaWMQlM0YOAm
Xa3YwMRgr8b1ZN1djYewrcPNB40w8fsS374wdzHVK/DJgAIOv6GOT/BtwabQnJJxu9b4Uhx/SyAA
4eQStTSzpGd1jP+2G9nss7NlUnyzulg/o1P4zlxFKiKSpssYeY3b2UcJXeXUymG41lNmpyXav65U
lR1W5ZD9GtiSTKYNO7LMJvL6yCA/McMhwl+iT2K59gX1udufCtWletfnefWZLZLUGIqo3MDSpQa7
IJY5jZ7PkHX8NqUQVJi5tuyHizvWNL780gzC7uz33pfVVvH5spHt8/h2dtC9FpYTlVL9Gt5GHLLX
LcyOXnut7JjChm9qJbu2zslw/P6KNF3zav7WwTP5+Dxo0nnnZ3X+4swJ8/8Rtx3bDu4smNMoYC17
zJg5Ubw5KONhkRfGowPVnOtOS7gwh+0lfoSo335HEH3oeL1LqCfSZxXcgqHiOGbZ7+Y9CJY3ORp+
vE6/rhI/PAmy5rphZxi5IJdmVWg5nYoPLmcxb7j3Rg4vh+sZuLhE3q0h+HcBtkbZ9WaQfZVjoqxm
iENb5fSWewUrCs8UnNPlhFLv1YUmucU+JD4xEstgCWLtBQ64Q9C0vFx0TPVUh5QsGwHMGQ1P6QfH
7/5TsA9a1BzoS+Tior8np3m0A3PsRByjbEQFLA0ogD78i6pbZZKMmE2wnKTvMKQam7yJaeVxgFLM
6HRKkQiZbE0mF9u3K0iiSOA4g7ODmXwHRuep6oJY3QV2nHiG+AWKMm97z3zhh/wE94263q6zT1gp
7xVryGkZI7zlIA6lfOdTOSq9Qh512yd9+mdoTVPZ06q+PQUN1aYRCBAoidRCoOWbD3z6lHLAXOkU
iALJUvOsMA0mW0kEVfKRLbHAqtrIh/TgmBUhFr6Is7TVGGb07kV868qbLZRi3i5hQL7wW8zfmmrs
PlZh+KIRE+BupqbElzNJYqCLh7lDFdg+KdS4crmP7hotlelrCzlEPmoKoWpzaQo61rESHCuazt2E
5ztCCPpyAtg4JXB9PA7KDI5NRTzA0yv8yTxBJrNKmBFG2IILtXSbHwqjLWvoKlkwCd9TTPqwHdD+
ObsmS/jOtxDB4oTczGM/at3rvKYAJ1ZzxP2TSta7pzVBX02/qZhZS2IqtIQmM8L1slPoX37EV0TT
Rb6hCo7RYs45j5CL0K0YhdbMxk0eBXjyTXiNRLdRA4QlVnXje0bIsfyBktY2aa7xV3VCorWBdTWO
iDdsRmAV7gUDgLLaYFIKmtF/puaBu8LuOXiUn/aHpzSmhAQguS8Wu8Q8y56KpQclTfeq8ldf5uuL
FrHZO5vcD18ypaD+ASlzBuk+GxIeg2zjcgjVNBx1eRFBmZGb2hHCcj+dBkMY/UK2TIRYtYnkhJjP
hcF4ROtkLol42B+7hU26+RwAIals+NxS3ZSSPSa8xlycHhaHokAloqY73TFs8WD1lhbxCIjWIL+R
e7Xzo4DC354OeRs1zJjQUv8EM4Yt3Ea5ZT7vvsBCV7P20daTOKt3DIGPcc5MG/WqaKVKD8QMXs+x
s5UH91t2VkT6WfJcPw7YSD/nci2jZzIJYlghWN1LQEJIIH1yEXRQD0QuwvoNl6ZS0u8sFsL9pCrP
xOCOsTr4ArYsXAnkwoG6YFjL53nkhCyu1YU4pfFj7u5nkkFVMjBqvIB8dyeDiXQCx77N+d95gUB8
HBBL3SNop0QRbFSIEY6LmhqdK/4FN1cM/EBx8cuOu9VDU62h1hZZRnW0x4shaDwgNaxb60PlPXuB
tfjG5YWhcNz6W/ocnnNI0+Sb8XykdACiSvfeWwZsJ1BuYRKewlz6LMKZxpSo0jgyxGrQUrMxToJm
/xqp2eC3JtSDUhfxDLTIl7oemPXOVwyhARm9zALha3VkBTah5X+F3xV+Ss7pz56cP7yjyu/hmz/F
6Mwl9fpZTYWReFsvHoopYpVOYR1J12q3Nov395p+dKaHq0+q95UJUB6WadJLrzCQ8eOQJuxLpLSA
o865WoaP2gtEAVgWzI+SSEWCn8fZT4tzmkPIsA2y9CmNhKMvwbuwhrVnam4ATZRcIMROp0v/cvOU
HdylpwHL3uO7bVi1VMqZzLWITzkEQbIpO/5XYHggLsjfcgSkeNxASvwik2dEyfYxYdORyjG5vjkd
Wbu3WS+f2yP5t3CaefADhVi2Fh7YsMZUHA17ucwSKhKel5squH7FFzhIs2HGAA693znihA7Tc82O
0HcyLcEcmE/MXA9GS7V4wsMRFq6XfPRHQNY1TC3r02X9TinsoKg/kjlhYxoWbY/Ha9/HgJBnU0oF
Qf3WFawZGJKLquLGrBqLZreQD7ECS1R0ffptDgWzuPmWN9PF0/vbjcSBVR7/eAIbmpp5GDfBLB5o
/aaTGBaJyD3pCBPjkEhJGrW8Z+rfYy/i6+3gvhjmX33M9AaF2mGEHC781Ia5p24V89YvIifyt/+5
/fmb1CVVGSaooZybTPGtKtptU96NmipWDXk82s7Y4H65ZtfQcBEdTPxgboWOzZTbtAZ/Y9aoB9+k
rQdkMnzjabhTqnc8aNMZEqdacevQyRpWKrSyeS9B9c0tXtU7pKFBCz4iU5Ec917A6x7JpQ5xlRI3
Mk/dL6y0gqcQscP5npV4Cljc8jDYauxlUanMk1HLrfjhNtwYogNLbv3fBdKvj6k75Nc+H6Mi2B2s
BbfCNGlCmw0rHJXuQBdC2luohgCreyIeMopWgJNBWExPkYJOUbK0tWAjfacIcUYh+PvbgXd55dIu
6g84w1w/HY6szUAE8S6aaGUa2iK6zSrlj4ztyvK7wQ++QA+MZ2LpBNdqOdF9/nMJmaAGDGI9QlLa
xV3MZtpOvsBXBZWmKPQmoS7Tc9JnMVJ7oaMMWPoO8hB5wTH1YDQWWdTc8Y2POAGYRkejdPKiwSTu
A3knJ9OyVIJHqh3MlPGYyBWOXqxm4UtR2pShno0O3joSRabNepRPZRG/xnyqq6OcR6I5QMv0DfaD
FSr7+P3un4px7KLcrqeDu6xSOq48uX+5fBGhxVO66OKuvSr7sA5MOKHrdXNxfZr99z6A09lxl1mQ
bGHKR+F8BQap/hkWKva+JWWsqGCciQRmzIbhVsBWJKBdHPRmSpRi5IQVxeA0btzyzgC+9uY6XaZa
Bk1z1h/31drRClX9KZHri6poRcgvWs4U70iPL+mKAXTnvjVv1NTqnuwt23XOXZ5ly0Sk4WJQuuGm
QtZdfkwFxWVKCZFqLhQ+aIxa/p5dN3amksPQuI67I/6PnHiV5NQ7/4LcfCHv5wAo7S8iX/jfX61l
54ZOw60Tv2uhyRhsrp8dC8UcDQo7weziiZFMuIC9xAcBog8ZAM+ZF14iilpuxjs5RU8/EQtuTKpk
AehYlDWaDMwYmlIkINhGqdFobzlrz9qRAXkRhPhxJh2/8PoYdjdlMB7apIw+4hTk9DnEJOd+hMHC
ccNF/MqZWEps9IjydKYv+Wcqw4VE/TsSaoos0BNmCjRYsy98zVQ1wiPwtVQd6nJHAQuQsXaQodp9
70CUEPjT/Ru0eSGv8639jva1VKhaHp1kNsuEl8v6sBlW0TM17589OvHSCrfFJOpSemFUBYaJGqyu
Nb5ZR8tzLt92cuOWJvGT2zYR9Pq/IzTgQiz481gz8ZJLyq2vASVspiV/1Av+E2kAcRrp+bZUJmkX
biEHVzSrEzLYMP07pNSy5iA89NtYwb9CYO/GgTBwWUQxGAQHLPA7LCoUKGGcIgBl0AEWwZL9U24N
tRoulnhNUA9UNIr0XA2ihkpSDOaaElk3QoiBy9/cycN2KP/33mR+4guoJ/XjQSildhHbYnMR0A1f
UL/oolzIdAXFoXHlN1DmXMH5ur4gSqT5GNgO/FNL+qiqAwHT25QbPTTA4MhP6IoviIIIjAlcga71
eT0+KmV9j+905h9zY/cIJ/1frgcp+R70TuSQ3iajjLBYkZ3VyYLP7DuWbdaBAaS8Do4Xuz+iyO/w
IP/OevJ+5nmEQuj6wYC4Xh+/NVUDWx/euf8omUhHPpnEShUzrkGaijk5ecCeiyfpNRIXjkLFHA5d
yv4b2q+3jWjp7u7p8Fxfe6LihuJDW0ulIHkzK7DYJ0s74UoSAciRwnLg/H9k3wgh4rnGnwPJsYgF
QFxjzoTw9xJjZRtPoz4mfpvcM+Gd+TTmNeDNM5BTEmiUjCtwxmuQjja2K4eYKUiZdcD7VVNh0nqv
FW7sRtE8k1TkMAXRLXa6xrZoTxTSVdgow75Deyr3d34t01WfrUQ0Xa5UriQjTLF0MFYGMU9S/5kw
J2rjU2rwIEdZNVaUC102c7h2oLdEluw4QW5LmhvwiL1qWlNarcHIIeFFvmQ5ixNhUk7tC5ShmrKF
dxMe6MPkL3Pd4qoCRsK1JO/ex8F9psD4aPno8YmzNxGvU0QBJjl1rXNPZ6XXxVa9qyWLdq7kPuFv
7RIxbwzy8BSSv3Ao/1w8Vs0rR0/GOKBr0K2Zwg1Pw6I4iXNrtiotwscej8QEFtJU4hnuPaZSIba8
JycWTm0+A8wc853bsP8RL3tRzpuFTamXw9bLtW35WyzGr5ctMZ52DpHSvZ8mQzZgAiOhhwROicus
tOmwvCkoVGSA3gcFOYg+P3V5GpC30iXZtLlIuqgZpR779xCiMKro6vn0H/sLegaZVYNFp+uxFRt9
0G8iWp5HabN5sUxKHEr68c+D5Cbys9oRjji+OYSJVq30+4m+qCgeHhTNnGLxbv2LX43rGVDCIxa2
/VPaxzKs3yoxMxWnGzQKoK2KD08ef6gpN8GpVUze405YP8gl24PLfHor43MJEewCWfQWgWeuYw/9
DcVFO6wNWvl8x5ffjVtJZijrtVo/+LTIDCyvx9V0QJAqdJSdaz9rSwHrfD4t+X2mPbLAzbqu0gA0
csNBhZpIWtz0brqqGDMSkBDF1+yuLnW4cu6hPPS15sjNzfdiX/qezMDXqUbt0ebJIaQP2ckz8ng7
5QdoMnAe+AYOSYymr+Gw2OANvZ3FzeRDFLBncvXboUrRSKhBCUQaOnzzeFwt6qKuxUb/DzglWvHO
WCWE/PYLgbXKNmYMxSuaz2QNvmzJtPa5t2IZzNT7LBSShblX6Wayh8+dkzVg1uLpq9c8ehFxEaXJ
4dTC6YryD41IDjFRmqFCkHLyizahLu6okx9r1/rDjCXmDRZIyswmk/0A6tJlXvM/sOGDdJG2NFIy
bJP1OrEkpvRfXxQk9xcJ/uhbnOk2/U1TeD7EOezQKt3xlA7N9jUmLI1PGWWZ7e7+7hKRDyoHmLJ6
L3QqBqXYw0SrHr69i+RYV6Ie43h3sw7T26SG81ziY0gS9YwPjF2B311CiQaC+P2wMZBnrV9P0HlP
BS3Edxv5iEbr6B0+l2zWIYQlEIgEhEKZheqfxSF17yQUh3tClNBi+Tbw82bDEXjUCge+ZKxapiCO
xzCQ8raL3fqtN66XZeOXPR+8+XjBtktXtcei9oXtpPJ2XiqjJNgcIS5d3UelglZ5DKtILPMimB+B
LD22dnl0ai6wt+9VoDqc0MEBXjZCQ3nnb5+o8EyH9+N/o3v7bRLhAj8aoaK3iVq6kMmuW4Koz4SV
tKTNdru4x3qnuwpCOLEspn5JxYNvjLyK55oW/zyZ2fQFiyJul/xzJ3EB5U9emNESz4+lgC79TS9u
A5M4cnp7ryxOdo5fmw45bZYerrj25dXoo3ddXk7kdL99yZ41LKOi4E7mduuuevhlMKWhai7v1fRN
+QJvmpLjJ2hgMz3KL7wOuNc7fbQ/cxBarG2OJ36+AR9BV4yegzxD74GS/l07q/pBxE9djDfYvydc
cdyDcAOuh84Z0Vgyr2tPQfMkl2eBUGRaBGHbh5xsm4ovop4MTzr4hvqm4P94MrN0TfmjUaRGOJ/S
tdxejpcCXr/aGuS7gXlibuNVQoIfkJSALqQQoe7Se+Vw2WCmQqgvBGjs+OjTMuEhVLe8jKsj3f3d
5HK3sogho+DQnSIfA42rjoqHRDzfCcq9YDryGnoP6QcYAe7Q2oFvQHzc+8+z0i+aWRVXKhMPwQLA
XlKydVKJBwNtg8v0JZhcQ+JmkQCL4585p8m2Xq23ieUSGZaq6JbKgxiGKwRnb63wklfVUO94sLsV
p1aDh9xYJonbCujyW9aOiRM5LJyLVv99YZgpM7CtqkVcVkTBDyGhV1dJFshHNHE8xXiRzNQ0Zdg3
UXdMvWy1twhcaT51l5AypolPe07HbHECPmnEj92QLlli9pCdxhEunYM5YKTMXyTkrCqBbTzqAELd
kbz+MP+sDkNeayE0wKH50NK6oMOFhi+9/Kw7lNMuqaODmPtJJE8CoZqp8pjcAs0i4ARkewXkDG62
aqkgahY5xj9ssFmx4cbDjdRer/yNxlxm6GsHlZ5XegGTB0EhAPnAaskjZzF80t1OD9z8FnS4Ld8I
ostKxSTmmE/piJTZpAzq//AvoW+xJ8yLVuKWWbkvFRl2QlW76LRvZuOkbd6iwWu8iBT2HxKXJbsx
IcYnpUtIYWQxRGQUC06iQtKDKlvxAEkBrk/9xkiC6xm5pUg2j9kGfNx+7gnZjrbPUInVjRXvg48d
nq9EmjcYDq2rg9uGEBVrdnhzpYuN3s14eFgf0Gzr6moeNvyHZju1tcS8GDogEUKxzq4CVwKVFPaM
7QRoJi8VpCTikMl6Jjcob9cfG9nx/FLLd2vulgct4QEVa3KxP+xc1jzdcJ0Kn7JTL5i6TnUdyzlM
67LY4VwoZFGczSvrALZIyrnOBZb3XBgaLKBQ9wcHptAOqxsVI0wNaDjoy/Y4Ao4yvheir2EFTuIe
cmQDPsnBuoEPxghhDQn3JZx3jpVwYGgQjfLF+X1I36Op+Ri2qA2mDMlhbix4zA6bWN+635c180ks
RpYB6tJxerZb2/Nmf89UpZalg4Q/6nIRlCU4WUrpkP345mjhuG4AbgG4VFqzwjTrnhyPoVRH9xrE
H7pdbDrPE5z5Ec8qnlAoJ6UY2rpHQksop7rCM4zkiPo/F/Chf1ISXoWBTJZ34wwgQ3+AO8G5BqsO
b3zOSoYG7Row8luDeqAkffTMpAzUUW1MDd+Ah3DWxDYpnH9qwW2dURRH5VtVbioXmkpoEnq3KQPI
aB8u3u+8jy+Mw3UF3I3IGkgTvdga/NBdruBJntQohGva6lr/iySjgzsA1fpawfQS3v/yeu0zUeNv
ooT9P2YsuyQQKuS/lTKeHe/WHVDkodtR+7yJLHuLtvlfncFIqYmOWPYEPjCGCOhiMsgDr3hC3Mlv
dnnPNH6kvqqRhM9QIMLZX/9cersaHaWxix87zK7LFe+rsj1XARxTbvdlvXTeiQhXpVQqzndRGMrD
bAWM9MlC72uYm5EnilJlAuNXfPwzPb/JCE/lxzJUrxEFqcXlzhE2+/eyA6d3F/I/I8jMUGDP7qyA
YbE3Po3uc6+XM7gMDwIsuNOK++hpPRUh6/riqUuLxZh1LObKsyTl0dGsWTHw6KSwRZ6W1CS6zP+S
aeoGz8fO7wdjSYNRGxS5b7JSLlTsN//9EFqKofCiIcF2CpbWmNCQsAMsS+umiFopS6ZtsmIo7E9B
Ddak2k9wRT/9gB0Y/P8vFPhmpmxnh3PLWDRptx8GerR0DoAM/qswHEx8CoVKxnfXACmnDuy+R9Ax
1Uvsm8NWMWYOcCwPBrIOsD15l1n0TsrB/IsX6PWbArDowOvk5KRJRmiD2vzwnJsyZ6sfhKgrwudt
qhgG2eVvRXxHUTbHUUFVvXUl0oENQRt/VY1rpd75hVUzh4PKLzag+QWVvO5S0BQ39gPA7KvCyvWs
XWTHx0x42H4IcU+Kz2gKuAW5j1DyihbWCCY4HA3GFoGrVAc2Ynz0Nd/2xUzatESKAayI0u+UKkuJ
5BzsmCKAEpvGEghFyh/6p0llbPImq7wlOh2Gyo/PhcgSUI4wUQq1NQwsn925E4woV9leQf4iDekI
97esp3KCpd+Wj9i7lwx9J0l2Mry3qDiNClUd43ef6ObDVnXt01Ju4DmnhUfeGmqSSEUKH83j9nJy
PMO1FEHUbuVRW8RiHZikpc/Mr7gixHEeDAJzs0gLYb9kO3uz8OqXdg5uSlRR7zjZg+m730auaFv2
ugzME9xwerd6tQyCERxXq5Hb00aJKklJgURAhpKedMJ/ab/JOg1sf7f7Acf7ZfmsD+8lW+oYJ0vH
RhwJE8MNL8QPIRS5e8rJR4vZM+y33wjrHYLWgS6IZo/3nx1aT/ZFbn0xtzGDzJvDR2lIoT3lu0XN
jDSrNxlUT3eAxmnw5B4dRMD4QLwtzQiICF1pOxK1xohLnulBrSFiiL+B2Wo29jUZkOBxH+AKa/k5
go01l6OKGyEDM5AqkYthOuQAlSop4BN4vNh7KKUXVW0uu3rWpEr9YdOuq2h6L6bOghoOB/K4GrIx
NGQiFsMhT4y/tAcr7ChNPpGz5smT5qcjsNWE615K+S/XqKVW1CMDV32gZy4rJJIl1O0TBGBEfujo
cATI1MCydZkeybqxluu4MsAcss9xMsYrHaXlwvaqb93rkk1Gi0ZzmnPjKiYva7uB4nZX6RkaA2bu
hU5HgJ3SuzVmV0rZMebtwm1NIeHH73nyZCzcqs000CjmCresldk2/KmZDVj5JlUqUSMdbl59kRMG
mhMqfP4lYE5s2zEkpUYyM5loEVxVL6y2drrnHhCC1+BuMGYMiYfTh48atLSmIIvgb7j5MmPp3s4e
Au8++CZj9x/HJ8ZdxsUiyAOELyqk12G+7Tb6OhSFnfEkRjImDr3glk+4OOe7lbmQ3IusExhm4W/c
LO+GHMzb9OxT9pEk/tRLWA8VB6rhEYpEM25A+GgHQB06d/fN1HVO1F+VWflFol2ML+f0KiN2fGep
HfFQUK0NVibYt9QcDsXgYINESR7HERf9th5LBTX8q/3aQ3NReZMv8SJMw8AYYlK+wF3XnZjiidvX
Ph3qVRFJzPetW566xuxQoBZizevI9B5kSR1cLmRA2nY9dJZ+viOgiJkiKyvJ14Go6KTlngM24dNC
QkR3UM1mL08a3fjNnb/3fAnZDWgPcZS7J6QQ6TCgZNUNyX8oau+lNKUsdVVr+9tiaRpLRu/BfbWr
yahCsvGi64ilmdA5LtljHgeZYh547stpbueqwnundFdQyLKsRhY0MOK+vN+/vAEDxXTDxKDnlMcO
SrNO97ZaOyy0JWwwIYvrvru2Dpz8rA9zpv04mCj4VYCOxMgC4CIfi2FCkafwLPklfg8luyNjTblH
CwmdBX5Yq0GcVRAng5iriNxfRX3B1JBwp+qTqNk5J1o+tsNIFjh0l8v2WkwmOw85VlFJxuINsU/t
oaedbdFmKb4q3lkSRDqpPWu9su2tO92sh3lDELJnJPVd6yKsSPzr0N6u4o2H6sDKdIIwxXWoNppf
Pqu1EpwzKdLM/D9N/VULWFFbA/46obuTSOJ5joKPrwsZlDuCl91UL0DteuBBwPAabKrHqkjnPlVH
Jw2eE2T0zQs+qNjXUX8CzgtigH4f00L7+jdpWX/IMjR29Q0RrWF50LhOgBc4P2pI9kmStlzMd5NS
pXzJ3864ai2kxZnMsimHjHcFlTe4q5dQ1bTDFJGZIpMt+OOHEQkDK2+8upXvMzZ5Ttx8brj97Q77
d5yUjGuckIxNjJF4W8a9FSPGimRuF/iV2t0DNBl2IwTDXBf/PjDXaICyrZw6yyk3Uym/V2bZEYj5
d+VxMStkA3RL0JuXJmHXs0jKTiYywMX2pP/0ysJQeyld8qVl3rd3TxJy7Ab47CwjCpbAnzGmuKQ0
wdX64aB/EXJubktlBO4omhra8HqtlX4yDgyTwHqPhkj50mSRYu/9eFwllcwOu5AdgKorCjAd5Okb
tDYaJ9COv/IPV0pqBawjNQtITLIViD8qaewf1NoDB9UTj8meDVkIJ2jHuZFMhbhwntJRYUQOGDyQ
xx/4t5L+0QpgTDMmZPVA9Y9OiGaQFVASNIhI6yxtl2YtHCGISLUbLmaZlOlZvDhJTgEmly9O79rp
zlIo/HWZI1mcIPb56e0Tba7sBLQ6BlwFJQ9XO7oghRNKTs1XSiGyBmJKiP9YC9LYcO0wwCYJLUij
3L1n2oaBAS07J0gzwGXW1x73fplpSwllVt8XH6HWI02QoiTv6eSrt0B9BGqxnLbgA30cqLjgZ0X3
iRq44h+u1M1qNmOlPeqN4jTp6dVM8GxR1rNHKrxOdvfpTcyagUjf+jgFuXjgK9iY4QVbNxhGoArl
kDexVCEq+OfP6kwAKRsTss+/zyZXFOy4QxYQjxGWdMx6urnaM7EjXXj49tOVlsLWO75IqKJKPoow
DHkrL07Ua893CeFzOrRbiDDvrJubGmC2bkxVYK8YWkMKy7GmK2GaiDBJet1RNYW9NI0uJPK4m98x
5G8m9No5XKnt2rkKkjgQn5s7IsWqftVRrGdwGVPxTijaYiabe8hKbJ3mKQZ/w03U7f+JcAVfSDmN
XIKMFT1Vx/UqAe9YiF+1K2NexKCA8VxtrdJCrFvh+pZfR4QMLGtbyzOzEBemOxXKUHg4p0uzOyVL
r1W9ZARgMZk6NCj5gOBHj9Hh7z/L8rCTQI9WLyHKY0sUauizEtYiEnC4weqL2USTyNW5DwfjUGlO
VNqMQJv1nxgCAxsvJmHMovx5ohMLv72ytFnlBVw5gPENGI71gFKPldnvEExcAO9gQhTtll0VCZl5
UX3ZtjB089Ek1kuJCUH/QcrFFkVJl8Vuc/a1R/f2AhfaPGqXnZdIjZau4mcjpP4oEtnSK48upGDB
EGsWJjLtAo4CW5I1jjFlDDSU6SeO4tTPtP7gdQaR0R+SK8ILc6Yjn00scF8mDwO8UqEgmbluuBau
InKpqrGijrFvCht4Ece3QjktD/ngKVjBWfu9Pa+4FYpg3jITepSuORb+8afBiTOQle+g+h4NMcxO
ZIgbYs9HOX4kQYds8ful6pujjhcvBYNmHieP6Ogc2XTfx6IL/6R3z8RyeMBQQrFWSBKYLvLEVRRi
0XbukvUnB88NPbjR8CGJYNhnNVR4A4xUy9t1h1FkAWku8iW0ppDxUeO1ig2ROyJKr+DFDQkFoB9/
RKtz3kfZlqjuyCo6qYdNT6QdZabT1Di7nRCNBDZbvJHa3bcq3+JxWAnWmpyUPVTChC2zBOaJzvbe
nVqwUEgH+hEt0XH3bqKSPgEyC4Pc/OwQ60voFB57ZZmK452nTAhyN9a2p4NPA/hnJnENWRTd8oKt
rWM4AOoLmz+sCaxpQQ5bsy8xDWT6zmewnYmRGEksB5ug5r5t09Sszv/hZc7BM2k4HbYRm4Zp2hYP
3Sx0jv1CL8y7yMLBZnOtlRwZfD1PIMrbVuNSbIWP848RUDHEuvsk9gLeOl4HsCMkn1pgG47OCK4L
nmH3X4RaMJaXSvE0Hc4zpach0m38HD0HYlGYab6A/zXc42ifzDqma03XbOWeKtDaMv7fe2gDWInl
iNgLJuwH+vWKWKW1UqHgcUkBmjmsgeSmETu5YHyAhicfV3SVuD0pyY48Q4Crmh865mIGda6FW/Dq
Sw73RLnXolhgWACp3dNeGxwJnUJHxRivmjxDYFEIOMpzAQvLCJgjovld8lRbQZt8SqnYpdkY1wSG
qOJa4MZqpT5rsLNSlNh6mvCbBxvSnUISTYbN1xuIGiM1PUxV2wmrKt1ZIM/fvTx+5XvJTjgfeXfy
W6jps2iAikoY3JIDrNYa5fZ2beJFwYOfcdMZzQ1whmiCZ03YSaa39IisO9DHiTraXIK3n2kAbNaZ
bLow9Yrh98LkRWU0M/clTZylM9mYWftujzmoGT+ge5RnyQSexjvMgJzD95rqyLvcEnGfZ4abppSM
m2r5+HQTdn3MFkWTq/8KODhmn1T4fJseuWdGCwlUC/UONRnhO1jMMGLnxja88oodhwl3lBhLGjrp
iwzksiojAglvoLg2Ece9Oqt7kDc8X8+HI858mgWq+44V43rNh+U/ZT7/OYfO1GNOSN+RWqQfjZMt
30Q1azepXePJ5AwtbHSP/5D/gkaolX6QKp1hjrBbg/bi55KFCbfS2qlLhaDSLcNGPhfH1HNUUBBD
qZSb1o8wztvy4bjxKO4ndl4zK1XTwEhO1QY6WuJ41vG3zf9aBy+eXXkCzuoh3IVo4NL0zoj3e/hO
NPlcw+4wmzuu0tJ7ckdccCGqUN2mdvVTh8tCUArYuggHAF1XDvLvY4AeBPFo5VdofnkS7ypZq9gl
6YUVyvdyrxeNX7mlZqUT7gHcen/G0Yuvy78WuYrpW3Ye6v/O64mvsSHDJCu3fXlJF/GY9u+jLip5
MMEst+gTCm5NEHcZTea4ze+HPqK234hAIMyO9K7ykz9+BxQ8NzIQUgkh0hPBS/ZtgMUFHWstEXAu
zMEbMY9pEV0mmijLnXSTaZ5OE7HMkjvQFj5fghiSBi8+TzSFbDs/i+HHnq7SWdK8pSOIFLxA7ZMU
vI/NVuWWxIh1REhjj42VdJBUMgkGTIn5w8mSO0JNfDmBPw480QbEXnZ78EHbvggcw7x3ooV44ENh
PjxqVIQP7S/b0KZ4lSvP7Cum+WASvazagBRk6a3Mrv+Nm8LFMXNemK6oxAGXE3Hw8EnY2vsNrYVk
1Jh9wj0kU6OXIqTLM3mNP4cf8WqcGNNB+sv8vZCcWW2thHVKI063k7bxODGRjdYDiZXn5GOTgvcI
0N5Ja0E0Y7ufKRcygnadtzIhTn5xyak9DdH4HlriR6RRmm8PR0NKHDpSJ4wqX6tXGY2B3vYfyqI3
Aw+C/zdHhTleTmDL1ApifQ9C+YqT5gm5C4e6KO6p7KmXmujX7W+LohbfxrekPsdmxu1eKO8tD2yB
4JWcZ/1NKlUrhYRD7mTE6d+yIOFuSPgEehmgLxBbhwtOcQq5ZBtfgv+rZ8i75QESuTF4tfb51g9p
Ejqm7v4LBCOJtriVWHmIwjkQ6/3QArhoeLXw2UHaPr/IcKzYts7fD3YmaF4hQdYuG7hS0j/Wtnwa
IRMjEe0KxVYTQPBvPP4hll4C7xASaASFvWRoayt9/oV6c+VjPQrG7Fr5jl18jK52C/R+wZDoJBeB
LPWVDpEZJjVkhD5cxW9uMVjD3q4S07Fg+BDF4DTV4PNKb2Hv+YXEuULo9NwoUAx5mgnGYQsbJPNu
9vUoDZiLMv74W8Kb1dNUb07WRDF2iLqXLjF6rKC2ftRwaAEeT+cYKWIpKALJimEff0czGIAueGzM
ThYlzeSgH7w6kL+esU9aihpa7Oe0eZS+iaFIIPwCY7EmZV9Kr+hBI02BEVhMOetu8L3UM8HNImCy
vqfEB+3VaayspVfHSTYZBFqxio4R7IDCNYYPIka34mFdv/4XSe0kCyEeH6W9+k6t76A9k13MTIAF
DLM3iee7nN3IWXOxWjGg78zKukIrKVgM2va6Xdsj4X3xLbvan8nLGKE31t9psoMRqPdo0AmYjFuJ
sRkRk0T9JzXwwy+1stSu0s/E1ACbihPoENWhuS8gdQIhRxXjFtYW67vLML6J/VD00bXAzj7ylx9N
w/sRs7A6KwSofE28GtO19M+detOJZdKyw4YIrHMvhCGaDcmzdtk6BhnCrMydMA5x033FhKk/ZlH7
wrlL5xmDz8VYNj109+C90XI6qe7Q6BpwJKzguygk1Z5SPCTOhZHUUT0R4TMRw0CA6Pjec+nk1Fwr
ouJ1TuZOiZieUorfT+XzvJeRCAiwDJZXu0G682lWuST3nRR3oEGddZlU+kM7M8hp44YIIgPizX1v
ty4o9O2xh4+RR+SNrzbIeUI2NfcmYGasmD5K8GOLGJHaujd1O+qcjCthBa2X5sdOoQ7SGw4tyuKA
+YPfyNodSGGXJNM9wi1CA0N9WkP3dm0r3aat8uiTkFRyoc1LmOjd82UbKd3LWx9s/CXOeWq/6aXN
asmqh7Yw9PyanB493FlmT0qyEofILd6PkgHh4RUAKzqRtHeEenvxScRUnh9z3fNdWqSSIPtvIwSy
9GOaqvvGqzUsAi6H82argHRFl+B7FEZaTa0z1wIHwQW2yeWuLCSu2oF+/+c2yHUfebQY2s7dhI6X
pa0nkHBNNo7xKrzG2Xie2KTz64fmFkxTGRx/wgP9OzdmWaUNibuRD4esCDHI3PbNhwn4iX7xab5o
U7kaUjqIoItqQAOVYTU1eFP+DUPR2WcMJdOlh9cB4s4aUFxlrnICh8qIBjDWUIfdS0eUMXltbh4w
R7C0xN/Hff7c9AU6/Xm4kTiRkny2M/0Utlq1Wl2awRB8tDh006mM6Id6IW4lC/TN5u0cXacoVLR0
+HMNv/VMrOw0qEJwptde8A8mkb1pK9SKcHGY+bvGu+Y4fF9NIkcFVxW79h7ecHJEJAahovy4hyIM
Hqyt9KXMuXlB1FLjHq5eKF/V533meFD1wifvgfT6eSY1Z+GGEiit4pRmtqtNrvc2r4S1USU8CjCT
hvcU7nRqe0m4hqdlgiolcPPnIoO65UxRPr/ahySQ//0V+KCHRJ58CiPzQil+8F5DWcXOw3rHWUAO
UfSZ7wGImpG3STOLBgvAa76aCMsjEbjjkDJVg8tcuJtEfGUBQTMteUQ09O6P/aDDi9dKaomjFpoB
na0EgndnUO7y/+5wBwrC+hXBd1JFltW3G+Cfd8OU6CQJt2qgaup9EKq0NoS1IgrNqUFchjwHCAry
55jRgEs5IpvleDdPiKeCLo+LOSbiEtC94zkMOkT3jx8THhmLypPsJSE7Le3hucFV505uAKz+CW5M
qq4y5pdF0jn+rBTJncQZd0+rtVyJEaqWwBB3P05ZCPtYe200TzKsyQ54lLKq5aWrOIJ3A+Z363A7
keSkOCxLpMRh9ExzOw44oYM/KDeae6/F/T5OULWH01q+edB6C4g4O7eRDA2JnqfcGHAsgi6wVI2F
k7O5cWYrxcVy52yCbsoZJBdZCWbFRbbUF3bHHKOPE9QJ4rLCfQnrMhcESb5KiV45PMYbTzSWJqUr
LrcuBL23Y7bdhGUzVad6ViiIG/l2mX5oTpSOxJtjZmVXzEVUpJA61c3T7j3INX9/cBzIcVsHTG29
7TyduyhyZaQ+qKr/Tnr+ro2IPRXQeVfbRJg2nZRZZagpY52D2yjJAWWNQxVILLgdYv9EAJF/K2SY
5q7KKNSIHOlahRlugTgOuaXcSTWYHyftj8pumtBc/HUtRB/aQeW9+Cd5Yo40Z/4W7v8PjYbDkp5h
jxX7FiEn82Q3LiREiZ5XfFGSd+VVL2vc0NnM0dwo/l9Y/3cLet4Qe8vPlwUxoHuO+CwIcXfRAqkZ
rLRxeLW8V6jI+2tv1BskbXvlAlZZmzQtPDucx3xzhLxP2/FumWagjgya0SthZ3gNxoopAtjkOOe/
c7B033ZERh3D1z7/6i6V/8yrh1/1ItNXk+6KUOJFxbxMeOxIx98BX/rUy4Vn2mSL0xMxZ8OWTaRy
Q6t6DFb0TJuKdsb+XDfDvJ1XzUqgE5lgSjY+B6+nfxgleAPbWdUjK0Rd/13TY8hrxLrBChQyk+q5
YpsDnXQrfncf6iZzNeT7lcwvZu2lHYCyj4uwctnYL2mfuWRRpLO/4nm3T0kmE9iywnfilCq/wGGy
1Qoundif2dTLq+Z1Tja0e9tBYNy9Q+pSQjVyq7Q+YQKNMtleb8bt6LTTcupCQtdgTKQjC2xhySvh
ZV5uajtk4yspZoMrlbZ0xFsC1q9P5WFpkmFk26NpQ/gDLJqux4/CzedJQSIZD79R8b45S6xBuvoz
X3Y625EKMmTTXkY4fh1Q8TZEjKO28WG5SKl6ycXRUPw8hkzaFZfyKUCsWMLImPjGPPCVqC6l2DqY
CBP+698hGkPZrQ9+kgZbzMLA5XsZGSUfRzaCA7SbI3iZUhrbiXNmOsafWlhMryfijVQHkZ+W6VA+
T4e2dswmSOXB86MUYTGS9XWcEijrazL3EukkNwNIGi7j5J7RaAiRGqrf/mP/zVhxuvm2oov6upIY
sAU0zmXsIvyIjfXkXdDK93qJBxFjQTMwOQoVYwRlpovU7hopi3mO5WRfKNQITksMeo7zxry/E11S
ReAaZrNm9GLkvXQZpuPnq5IVnSlDl2B9iVwWInpP92+hvh8vMwo/TXg9voA7ZxSBr5k3rc7DGBPJ
drEQ8aS3JRHJ/g30ImWSu2e0mR3UEjDLGTPRbYFFW0eUMyJaUYkH2X9wBEKNndSunGC4hv9ZUVKr
+hWYMVaPGianzaoCcJZ3fzS91KM1erPKT1IKj8GQRjHbXxUNG+z5MlmqPNCtnBLxWrAPiKQL8q+L
6hq6j1spDYWO2ojAzHsJ6dWM/BdvDLVclSJIQvAV5xMwmYEIGFHeL79iU0llZ1LkeO2Cet2E1Ohx
2hm/JbawQTz9SCF/uEXVClx/FgpKlUc75x+2U5YWabCmSuV0ghRqBFUGVR5baMC7E7pUei0npZlz
M1jc41EUzSn8aBr+bpYpbBCFJLU2O1qisxd5Di3f+M6L1zzBpQ5iujWqzpeUwYF3h9Rve+5LQof8
jj3crrJU6MEKfA90U3wbLCJU4J8OBtCDqrXe45YrzjwsXBf4vvJAjGraabC2wT41HmaELE3U4WQj
TGPH5HpaYwEcs1ThtyG14DcSxvTKHEvDUCLlE6oKqDb3eWJNf52X9/ZZRBrHWFhp+iYjhSR0daSO
8txnfADvIvDCpik0PsT97TPC86Z1PLMI/vecuFSKabAW2WDQg7VYevtEFRF94Vfh+6xQ/WOazKrz
AEaDrdC26+NLJXI5bCMTLzDS9XlVnqyoaSkmJQsrAPXRV+QjKH99OSJpNncKbq1d/cVEr4sdx7Ad
dy7bzUHqVjpPwdEHgOdEQ9HTvDraj0Yc/LhbOjkjCIL03FNfmYnCfurenvdJ4u3W/IxxTD198voN
NTciXGBI38DGGBuiXzahba/G5IqME4l0gDPjxLcSUeF6nqMT4yHSUFjTCfI0iIdewoWBojdH0ZlA
uFz0fj+N7vaflJAgCA36NiBi6qJFX/dkwjbGDbIpjzzP6E2oLBGnATIZrymPS3teIDoVZau65q5+
qJjAmjNIaeTzW9/MAROO74gQP1ul5SvWMc/E/a1N/CuhXoQK7WBxhmnJWBJEHKlc8+0tSp0sGG8d
zN/VAMfjn7VBRupBdmFWCZ0oHyZULY8WZt1mljOOKS+BSy1IxWpsgbGLzqebsotXwVtkN5j8ZDo3
Np03vXbESZfUdBdqc/bnkooNcTGQ5ug7SBRAd3MISZijpBH429NQYXeYadWSAOnuH8KvE0zcdx1W
UnsLNeS8QZZ92vCPxeCNHefEqu+/H9j292ZYDpbKQs6UkYwYQ524mGbp5YOWuDF2AKWPIowux5vb
JGKzugKh9ZsATx3Th6iEnOg6/JLaaYVJc8JSjLoqSJy3L8ja6aKanwlbCs2QZFMV5i78vEXoGJkC
ImpIgv2+22BT7WNjhViUN5nf0hcJ1UXfV/FtH94pvPuxoVEwpUkYbVw7iSMUzxY+R677pq5riuEz
dWz084VnYxHvYPf14hDDmx9GBt03X5KzeCk9oyQwZvxK4JWBxRXI41u21Mn7jPgGZn6kPdGY3vex
8UqBD3Q3x6dUiJcSdq3vaufrIuw8ehA4jdZiksHfr6Lmb/SoCKrwzX9HWr7eFSAEtC2lAM9M9R48
ezuYyG5HaHOLL9KuIxW8qn9EBi6o7PMpO2cY2skaTtU60w6A/PjKxMkF6vm8NnBKroAACLEyc9C0
bF7ldriuDxAHeb+WOpC4ma0kyyPS2djGXON9DjJh7zJOn03agP+X8U2fI0xdFN+5V16juJ9EWbxw
qFZySoWWLPRloD207+HDO6+IVkNDexGGAi+rtXIakafBYBzyMdTB8MTPTvfx2P9vuj0YoZM8/4Z4
WfNdUhQK+G/7P5oh+rwIHv3gYb/68sLlROjNU4Jg7TweOacQY3AQ3jkODOc0vVqkMbZwukMzSBAW
/+hk2xTqoA1GT6gscxE/p0OLfeUSudvn9/Xx+BoD4PEwT3Nm1Zzl7X0Sejga6gRy/5YtOpRPhagQ
qO+bvFZhAHR1oKl088GzTkX9qppMVGkLQqSqV+EC9a6tCDWar88qVTe+IuTGesfEMIx2QGhZE1M0
LSgBih2YlUeHT6Hvf80K8+PwyeO2ol4zeCqa8OQIeRPZzxnhZ+93XFXhDEY8WggSdvlKiPryKrLo
1w2vpazy7hmYiT6hIZYFReCAajSLTzg3s1m8V7RCRUx45rgyx+scWL31gXAYUHt8hCxiyZpf499D
9Ev6BPhZccBrlV3/zd9guAR9eo1076JCYWo6e5FMcCmDnv4WTCUt7osGYTPm1Y+GpGPiGfc5xA2C
ROTn7SIpFMmLIateU3NfsaX/enf4fK8hs9SMy/NbX+SRgrpmVSRBtOaqr/9e02wm6fAPNIwUgsom
srTK05H+HPqwqdEU98lb38XKfFpds0pinpCYdMPfmogMXUcU50RohPGIhX1/Za7XcAj/r0tJCKMc
bpxKUFUVQvY+h9jp/q9k2qAH6/iU9Xu+KPT6Z7LWIEhF0Wdzn2lzZRCqXEZQvUrQqTmwWh6ebNg0
pWh/VYBRegN/Y3PQP/ekGKJQwgS3b2QCrlckmVFhkw+WBrjXaoXZS3ssvdTt1yFRn8geepHGKI6s
Xt45HMor/FNqirlaKW51AzPVzmdimp/vPVZ0KsaNb+KZftuOsNodOd++HxVZiN3cRBE3gLNWtcSt
rf2c50osUlk5Da5RuHT+PGdsdM/BjEsnSTNTEX3/gdB89Juc4mzCD0tIacXtxzNGPzg5DFNOBXPJ
t7KzDfnfeLj9KkWP38trY4NvVMPvzeIZrt1ePXZ07X+hNVWWkCqXGJFAkED/QSB3QRIY5LmGplBZ
qFygRch1M85tBj+w/6Z670nZJuIZ/+VNfb/QwXWPK3R+yvPbM6lFeePHix607KaOf+zuVspEHOBt
AxAJRCBdqKcwD2s6Xx6iJd2ByJu5xr4UC9PhxTQ0XHK1HolCIfokuJQ1v1vWM3JHAJcXAv5599Iu
uH3mpMoW9/v0IW2/dYJo9cTbDayA2OqxASqOx2+mtGeY6/Hha9vE1Bsblo4Fb1hGARiIGry6Mh59
qNb8cxWJ5+kY41sb7YXxClxC8+GgJPT/Uyi1ZUfudA0cXpZUI7q3qyrEVzuOKcboogmvOlVZur43
z1gUWUCSCwJFkVjsAsEkfrKz+RcSNVJgjg6mhdhra1wo5Dwnwpu1C/V1GQL8bj7Jj9iVqoB6PPI/
CZBygrpO6tyUcaApvN422Krpjw4T1TSDiaIrFEt7TUCkD8DP7rO9v6nR1ylqeH+wgmTra7EMHajs
NWQn/QIYZnukVmIdbnaFvOiLr4IQfZIwSz8pqS6CWvcuJnxPDaIYldnowCXuM2ZSODTMp4cI/3zX
KrYbZPwZwSrA3e/TEVcyYdXBl5Z/P5dN6IMKH7YNkmZdK+44BCAOliuSFO2AVxlk3tG5WDajv4c0
5vI0qUPqGRx80rT1R0T6GI159dQC1hRPoI/6zSBFFvIjV6emO9kIKVKVrQRkvH1NpY23ZoxpCBI1
dXlhMCx1cz6DZTNrickfnntTnePSLSjxbkWUQW35i4kARE+D+dK3T84yRXS3XTgCbQspf29F1wao
EfSbKHkVCPTDhswIMAbjz+qYvIWkapxhOa6SRDko/ONXWDde7rXqXlqjpmqX9zbbm80zUQdk988F
mB+218YdVLsOdMN5sVD1rbhE+c9joRguefQoBcfNhfqoJrDX+G/Q7JTgolOCDuKtpHcnze9Hr8es
+bl9bYtWl8Ic+pFvm98I31Pu5+d+sZA5QDmqJiwCls+MrUSqPeWcTmTXNJ3vPR/V0y6jQJPO0Bbg
ezmh7YiXkrRenvFnDQ5fgthHjbc1dBvGfEX4oqtJn7GIgQlpkX9+EgRQ2JSW5WvjNJ1NMW2VOJ81
7K/4emISFT9Gjuh9SskDfioTf/xaSf3m4N3BUUeKelTREdYfMV4kkPKXSw/9+CLNFxrTHqLLxY7m
nyJNC+2NY8FO39qOiIxBI5X/rD6tWI2ejfiRbmaPUaRPllCSo9uAZdbysU/K79s6RFndYfWyGYTS
Pv2BwEVTC1i2KHO2/d5NHQtHaF6zBojxgFhHLxlHN+5qjZkBeZpNUWha9cFZ5bF7pgmSWUhUCZiI
kjNL+e7VE8Vp9Ay70EMhWOXFsrlwnb2VAyEa4HyrD2KVWpJfazTa/6gn5JNKTZqMYMEATWs9pPbK
SydCFdGJ/QToIxU8w8xplLxmMKfVF0Sdj87QBSXd6v0KQZ7QFDQjtMz0P5YOS7ScjrgY+CRvxgxT
tOjHR5Mrl6QC/8METWM2vnvrqJ4GKFW003T56NR+V1MhOKCKt7iYiyHGOs6k+2HueZJqWL7loTYr
RvUTsynVo9TVbORTmeAtaYWiNpKL0nVH6DLfeUp0y9giFmAL7IG/2bxuiuPtnWJZt7X20EJZCxj3
fZ9Pd6LLVWCr7zCEAFDwVITBfIhclop4OmZzLNnH9RlDjvFnZIvbxLj99Y2pRUhAzJzlKucFx/Dy
O9109huqRGw5kqmFVU/EoAzqSm0Vc8JBy62ZCh35wwYcmJ3z9OHBpmDHLDo0C14r7vqL+0//o/8b
Wa+jZDx2tRgUMJ/DJWQDN0A4c9N4mL3fz++FV6e+4m8d9cw+Sh8BeDJsuVYk3CIGfRmIp45EqBhk
c+uINc6YKEWOLnBvPlLj/61sWFL6jXda5rxTSKB4Zvi+iShwQBzaFn5o4JIpoxGVkATvyej1A1/g
Ex5p7fLd6wpBAfpc7PubXGKQNGIAgKjeUFbRjQdqesefMTrzZXIEPMYpezWV6hkCOEtH7abL/ol4
47s7TupVTQyu7ACi0JcxWja3junR/WfJ4qCIKEIpR+uErgI6kaylfExLHPGrDF8yl1MfXSfZ6YkH
e3BY6CHUn3V98wSgDKXk2gTZNFpPNLjWavnYOkSVx991GWdUzdvHNoPSH0K+0AWYH7OifzQGpm3K
teqox+8Ps0hmoiUYjgNcoOXysaAv5RmTzk7aoF2GGUqycAA5RsiQJ9mdmXbuUigdoxbyWll4Vco3
9MTZmUeqIwhK+ODvZ13WpxC7WMdqmeO3q/iJS5konnkGhIbm84fRxiLcNAaYhZIVLG4yOnXvVXUJ
urMhqZjA6ingasFo0UyRhcRV/N+JL9X390FTPAG0Rh87Aok6MvivVKN/3GAfzMXr/SxXtnhptxDX
5ui+2ddAI1BOc5ph7/oZX257WQcScFGG07ILWdIaq+uJPsYK7I1JmIpMeNHj/dPH/rNIASJoh31l
zMya9ve6QI7Z9si8ppNTvtzKqNj3VJBWMOdM/zMgUIIYG9BjtChWCb7kZpkZnlLA1mk63cDoQcpG
NwRTtZGD/cDwIKUedbDW62tm0ABfa0B63JW4MpQ8xg565UIOmi3jiK5za2klDR4Jo1gFMEMolrjx
iQW5/AUOFl/9VO5yUh9GjlOxxcJHaOF0ynNRmAhrk2+l9G8SbT3upv3PXi+Gq9Cm8Q+apsRxUbQA
QjDso5yE9aCzhmTCgF+CDCjXucxFYwXYjyJ8NdtTqChzQAsUwgo5ACCI71VxqZ4dDOxNv340cQ+w
Wf7KrWW2kqCrrkGLEeWPX200EQX7oINlbaIBTbcWWD85XKipkeifIEfGpuOXXWja0ZjiSKnOZdNv
LBAUZcnlhQbr8iHa2yb/msHxjPMH7Z614rY3Y9SaHsOGQyEargtHFjPvuGAio4/XBX3qaYAGvyHj
YKs2EapBDPSgycDXdmY+p2fA3GAs81RjP0yur/kvpB4ITIxzThWdSMhIfBme2T99msd00gw3FD5Q
6MDEJVG10PWasUff8Mq5n6aS4nxo0z5FVpnsTmNh7iEwr6Rm7tBYNoCYrzYrIxlqPCxVHV3cAybz
EViiOOffOkt3LbZU7MZRyE3JgtjeuP0mkifqPv/Q6y6ccokSgP5lwFSCVdFfotAE/7vxfSoNNpwD
KktpXgoSMeT2aUddAOEbF7WCtA4VYlWhZY1asVahQwpP7uvX/tI1Sjm/EWhCbSzEexPickVKTsy7
zpuR6FQopy0UlcmONYrJI/AIm+Gjqv1IScR2kf8sTyLwJ+JKwy5Yhe4hWcTq0RlLE5cb1up5UYja
gRCqgcEVH3Ky+YsBhiWcs+DkjkG+g+QbX9tJHtxq8il/Jsm0T6Wdut+zNMmMxLhixZ7f2Sw8jx+n
u+zLfb72BjWmVCDDzvKC5bjREJF4I34JwM9Zcr2cRzkd6I01FM3RgMks3XBCnvARugar0JRMcfir
fMD4Jnlnz0WeI3AMdrOKm50sjBLT0klMy99ULXSKcFBwrDOI2m1IyfEq/fK1vpNBm5+sD7X5kjf/
eawzmJUlYf04JwiWNh572Bcu+L/b4PQfQO6Up5nYIleOxW97dE6XF0vHrTMWSNkImFS2nUulO6/r
V3aQ4vnCtHB+aP+CDP+mVq1Vylo5ag7jKakl2RBBqCBAlrCAwk/47g6zKbxDzPBxKyY4tcxvBj8a
VcWJQRbdqPsOABMW1fPh0ptqTIlpQSq0tvxLDLoPQbFIsLjn0DfLdbd4erQb8zJ3qLI2fRL3EnNQ
R3ha9F3cbtOCyp44LoRppUj6hzCR+xgs5EY0snjUPDtGm6BAO2F7H2NCgGk7IzuasdL3xOw6SqF6
HyUu+7KxPB8kflNKJuIgL9/ToW24GP85T7l4Qn95DjDySc7oNBRSJxtgMyj04gJuu+jrL+/+rM0N
NYVAQ0x+2ZilWNOryt4Jnzk5GICOZQKNb3lIjjLGj7uMZ3Jq7Bqz4eJU8rXqiAK/bLjwwKgweraT
zt/mViCBsUFQ28W2y21DMvPaV2PneZ/DDzAu/ASUV5BEP7kYVZmy85gtdz+gEc8hQ/BF2qkDOwdF
OglNPk5/YWnsbegqyWO7Pr27fNhfji5B/JGw8mu0hbjS1Saadpk1qvoTONMQk45rBO08jSKPvfRa
SO7Frll0VcTvApPfMfB6Db5/M5nFvmFFq8tMKYmBeoSQJp2pGBqcKvvO4F6tNj2R1OB7kmFoMqRT
O1yImbzYrF5UyVfzbTq6HpgD6srEbcSSuvVWVG5PRDE7iqzt9JesR7UogXNchUStI7HOssr3sLca
mNpkmldnki6GbFuKcMLZBF+xD4+wOe+dC1DxZw5I6P6Kv7x8ZkSC61u07vRefyJy+vvY6a3Ij8Wd
8yJCtVQhL/ciauER2Cp//6pQNDJt45oai6uO5PHxCSxt5pIwvXuq7yqAlEc1Op0zrCDx4irGNkNb
jPqRzBAtN5PVYnuB6RnwjRUN9f5H66IbC3agOIDbO9iCq+FVCGTZVJUwngLrDj7dfCYLltVCMLsP
FFRUiFB9Ei1GJsdHeo2BJS/X5d5BiSZ300urx1OBcQtOvFXFcvvIZEIt23mIP6psMO+ImMUHJt6U
mT/hO98wt8EfTyLBhLV0zntNVC5CrzqhACRBHVgDTbaHMItUFmjsiy2clzluiuHQ9zL6F2TwQWjf
Lc4yDb0PT+5Ko1ChkAJEGlQGbUJfWxzcTC/9Z3enljLwCSVqzX34cuDZLh+yQoyuywF7tGV6JxI9
j0ah64CaYglwV4xkuIuv6SYLKGR9cT4Xok7qP81FIGyCgNst4SyB+myxNF7hdbFQqjuuVlkHHDBy
+9hXGz+1pSQZtCzJO4tGixHseqo2+a+oRigjjBwTesGv8fbhlx5fX/kuVWuJt7DHvSVJljKGWDVd
IKdYVobkZMZsOuKxOtdcPQYrg1/+9n/uGERN6yplmpa/2gpwbvay0D0vAjWt+wqAN1UAU5zSh/+a
Z0ClmeOLb2m/IMiVpJy8hQZZ6ezW11S1gSyDnKvL0CjyDshOTKjwtYWLro1YUXQXKz2fZ/9ZTdco
eA3mVYN2ioHvdrxzeCPRY0E40KdXxQGfMyjl/hpxcuGK4aRtOqi4gM1aIAdv+MBrnvlhhEg4IFH/
EGLUYPgknKky313dknJWzwQsiPqPCKlI0CgIKDYbA6XQolRgKE1BVXymDoAJQVKN3CCsfzWaiYMY
WHHeJ9zJOmWf40so/vuKK2W4GipwPcGrJ/okRNNO2P34fF9LaA/9rvN2ZJlKxPrGB7ezA56yAIrR
eAnTUIjZM0YTDsXHn21OqulAgOE7BH9lF/QJLIuZy76HI+9tYjB9xWNQrZYp0BuPBWB9J1gUXjpj
CHQVedaF+1mUZRWPqDxul3ISdc3xehGX0RBclRMJPMtRCgqJwI8yNBnFSpz9Pw1n9qBHC02Gh+P2
wbv9SYCEw3wf2aucVy9YL1r8+7ZhYxa6Qml9UcvRWNNXdGWvfqsJ1s3Cvkki0JFr5Wask6gedWnA
vyLmt4bOaxoTkjPe1tQp4suxFCaMj8wAFbJcRjnjTnadSxynuY+fji8YBF3SjoDbTycsFJacZHhy
SvNBt+MOrZckRXamFfupurCeTlCM8/NQq1tbH1dejGDfeJokkQJt5xeJuyH8Ix+cJWjriFk5x0QW
yBy5F8tMpCoPD+eevRraOdIMfT+gomrw2XVmpOXd3fbG6xqHyjdq6+G/YdzgMrDQTUzvJ65QAc9s
kimKku4yvGAo2SP1NQXfXZPV74iSUYZVyUgKACtV/d+Lu0qpyv4uBTnflYqiLxFBR5D4sHFSxyE8
GyT+lDV7Y0fflvnGUqP7Cdu6L46gMHIUnngAOUK8TcVRFKI3OlayKfbK3oX5PDnswUsbsWEqvBaq
ld5nTi8kkKyryWI0fmSE0Ck9Uw1de87n+vNleG+Vl4COJsbvGqodYI0EcII28r2QE5EnNFJeaoFj
45O2xK6S6JbKG91ptjCndddptG/iObQiwjijyUL37f7B9RaFwTfmLpXa4yoxLfsP8TBFvU9rrt7i
AfUlR66qmWvrZSZ2NFaL3xGbPZOme1EzgTrUpUusACMef1yb1iE0xQWXdb9IGHxhoPGa/Y+H82oW
aeP7WWCuGM8d3X1UXiLmdnrEoQtdr6R933C1+VlDpaIUnNa97fbvtYp99q+fIUV5og+w464ZmHkJ
Psrz4hL1urv9ZvlTjf0oLKJbHQNIr6v/Ddijfm2W7yA1p3rpz8hohBtC/N3RtSgriLu6yK4h0gGm
rCo3x8Y5CHw96KMgnBF4qkUyXdyEzzcpTev/wpIq6WNsETvxoybmanfZLbMDOUNJLFajyWEPNDXs
YtZViaW1tvYEzHfE2pldFvK6H98FwXwF5P8d4q0VtAID0qu8RR/lpZtgELzcMSptxNVkjdkeyaRN
5ohxIgax9+VrmjCihYbWmOpUwU+aK89hHRM606++RCvVggHFqW+7MxRVOpM29+Axb7xI9bI385Ww
ELJWayAyoAgDMkosMYy/tLB/8BpKsTAa31yHw0pbDeL2NCZatWvbF654RBr99r2w6Zra3fLJ2EsS
34hf9I/Ei5lTlLvf0sgoWDYAJbIFpxR7hE1xDQJ37rha0unuRQEUwgg+egWiKHDPdiR6V6Y0I4Ht
kQvBVzwni/WR2dIEP1NdB85VkIC+rJjm0xoZY9abxhtAyawS2fI7NZIhUwn6YT3Wo2iAbEhEgkp/
SeLM7EWEs4ddHshT1WRJ374uWO6gSKhcBnPIKzEBGsMJ/Tktqq0E6z2MITSjSJyKKWSBEsB2Qs9N
DlotB2Brfk2P0EaX808DPbezSPyvu5DIlQXephOo2/foV1vmBCOiOt53+zxoWayiVNzSdRlU/AJ/
i7mp+4EKR+XPJxecxFOZwlxhSG6w6OvObyhjVcqggunNiSg3u+1BT2RViB18RM8S9o9/5oVpTf6i
H/e/XtjowMiG+t7b1YaFcpapzbG0h3+fkEuFOl5SRS+jYwiQCR08QcidpbrQVV067QwIMdOe1i/b
LT0uMy8xaOFiW22QQs2lJyfC/P0E4CL3Xs/MZPJDHQ36MRzysQYKb/wP8z3btWENyTKkMzJ1/0Zi
vIixmAMnIouBXQF37wQ7Ejv4QcEBb8wF/EF17JRhrjPYNkr20TpZxlTmA/Y97rWCQDf3qWIdOLvu
fQibjNW5ga46pEsCbfPuOpmBlHRXY2kxeisideX7ckG9gTP7hBhC/zyXaXkG98YCssZQjw3SqI6Z
c17ZE6mRlP/sdMmBArotQpfXAuhzz4MeC6DRHGneSnVdE6Y7ZyYuYEfRbEASXDt0fWB2UiW5Hseo
W1e2LMUksSrT0eV30WBu0/ECO2Z5Ct0ZtXcFVaE2TBabJgbnbicqxKtBsGemEHnc80k7wk9mdAQi
NZA1xzNtgpkrMegNPQkS2T8AeWLIIrCwh5H/+aBRAB2s36whC2Uv6puvBECoSIE0mGg88llBtpEB
96pow9XrCH7SSPCkaaLL+9aBo8an3K6i+/aqYA5zxQGgDQb//z7vxoukbFAUGTPY2f6hQgTMCcTK
jTAAMAvXE3YAdKt8pIYAwkz7KhGcraJcIGJYqVx16BI1uSaBHgGWa7RXezEXdw4sxDBJyus+iC0Q
qWdZws+/iAewbe2ogNQ6RDCX+feej28kniZ3J1uxfworSLckThjCAxbqWVgxY4lwMvPjuCmbuCtG
zUecTV1b6M19tKJCugnKNa+QAtFgVqqTBDeOMkwXuXqOgqmaKHSxMowzRFBoTkFz9IXQwA8Sluo3
SQ81m/BjGrlUFK+IK0A2rxIPpseMlv+Bm/Jac8ee63XyW0QwSmGsYugYFKniImUa4skWJiQESAUY
aECLhMcKVhYHFo3kPrVDXkHIE/1vUwHu9zT+bbm4intG3dFCLoWNRPRVoU9J/Iu68l3jm5E3ToKi
Mm3JXXh8l5gpTPlLM0V5naPltLP8pvFOdpw4tyTuCCsmxKNzRe5WrC8kP9oQgBwNU2fCWdQwrRam
mzvYuzdPEjk6PImC0veKoChWIYl/hGcBuIJhizCuDDBHKc0nDrFE5AsCdTlH7l1TI7rFa078/mLQ
V1gyRKB6TwDRIztUfbE3zoVSH59Sm/J63LemMM44JBTXfaLSirZM6SvxRlaLIBa0LHZGtS+wojZM
8WSJECVBD7O/35S0ufkBEnWtVEQpSyfxA3A+bwQXYw/ppzJExt1j6DuAWdpjCau3XogYDbu+IV3t
NCoyHPZZtfxoclUgWl8uEW/jONqPo3adNEdCPfVHlVcydJbJ4Zb3FtCWpWPx+Tahq0ZCSBXuk3fb
iTJkRaIsuVJS2OvWOVfSbz8NHloamW2NkTBugHKG91pc0hAz+4PvOb5ca1YGOgyZKGKtScLONQRu
saSKVu1djP8vklvpKfm8WilFIla8D2401u7C5/q3K/T+gwFXAxIbVGUIsbN+nIwMybKslIwzqGwd
h6I1zZ/2CqLWuMw6eFHpObDNXIzP60buhDPj7zc5312zVnyIn6jPnX59+s0h6YmlhSYMPQ9giLR8
NlKv3Ky6HL+cqQN0kWdL71r4FM5chUhKi8HJkgwhfT/MCGAdzSgz1zO/iWRgcjO6yjZEZjm7S0mh
x2oyxrOqA9CJ7A5Zhe+Uc6oz7Unzvy3HhlIrsiTfa9H8hATxGMYfX5XyjH/jnQbNlsRA1yrARj3W
s/Ht21m/r5h9i7bxiSPYywBnvYUDfmyyfbh2o6orHUxX3wgW2UtgluulfaLSZOfRXo5E2qIwZNLz
c//yMHfjazE3e5IFoPS8UfYxBf+jNf7IHedYayEODDgRBBTaZjeMWa0d98kmg1/nqk7XAzlZ4QiI
aTIOwhsFQssylp8YdML4ufHRAOKGZSmTHa2fGYRhPY1OJX3Hh4LP7rYsWskWHErg29yAg8jLgY50
9X4jAq/jIfxiHJ/Lq28uQpRI0KMnSzx8rTXB54C/smf9ntp/m9ANjQ/5OhNwppwd1U27jWEBcsjO
RbD4L7Q1UB6MnbbENgEKMKj2ckga/pXwJSeGQAjznzjSYSLG1rm3sNvGUGeEOeX0MV47Dt2B17Hh
xqWtd6h5iPP9a7pr+nSzS4Ss6gU8e+I8oy3+9dPF1gqchovfBQkZRLpV62VF2mSdXt/PZjiOIna4
LYX+rE/EuQjB0Q3scQvJM+noy5b2RRE8DwYxg5SHafg6oO16YPS3dxz3glhDSpShv+OIsRSIIVE7
igLGvm52V3D0mzw6AYD/5a+5CWqmtCApwxbUu5uJOG2aGYffZAY7DKuLvi2Ziwk7sOxd9NQX4nRE
KQ19+0gZbJpie4X7Qdq+x4p2UTCv+lAgqEKPhadeS7xyWfMiaoyXXxpv2OKS90qkr0qd70//8tag
0IuIXlWiE30JTQIIHc9QNCdhf6Nh+2Nror2yPbi3OeDE7VUnH0G9sO9J9RsRtF/ic+334Ii3KT6p
YhPJ8RBEeYk/Y1peePE869XUmpWYjtptZRU4wVobVH1OexvWg4y0m8Pu6UZZdAre8cCoAFamV4dT
6mANK4Ylj0P7mZImA+NXWhptuBTG2DGXEdg+00QeQ4xPaYk81IJ2OwWnD6j0emQJSuQU/b47g0BB
2UmexyMOfFrP2Dydclco87V93Y6OI9p45IEM8LZQjGg9vrBBVfj3ptl+LAqIGvVSX8xqqMLN4P2y
o7ZC1lqmLakBarwu9EasgxpKd5P3XjZearT2WU2eBUKO5VQc2QeX7PWUN/W6ZlJCD6VLkLGr7HKZ
e2f3SxwFYdQW+33fYt+XKY3FD92PmKAE5ccynJj17yZhwj3FQphr92+wsT5lRKttZqidM9Yf4txc
0rQJsPSLtFGa4i1HKr3KMM2oR5liofWJtsS6PhfOEYF0lftUfgKcoXaNWBoIAsHqwNVUXnn5qlfg
8fLgtN4qojq4ihpnopZR4w+v2d7XgH5P0pn3xW+GXYMBr6lSZEig0XnNcF8yX5QKw5yqDrnphu00
Azh/zZ7/RgmlGZiU6oMcPsFvv7uVgY/41JkKXkRT6LhN5QiLm/rWpucYRa9Imb3uo/maoPEw3MW9
ZvFGpm3Is4W7eh8NShppGUOUPlRcdOoTF4T4ZQdtC6dtdr/EWw3Qv61sUHwJW/YtPN+Kul86k+h5
YP0HM5S1WoY/cgCjA8rrgNjUxiFQKdRdvivrBDJFKqm/cnEXVjMc80CgKre54ru4g9YcGlEd+UaD
L8iLL9+TTZdtGjlnRN7NpeaShtKs2Cv9Hw5NT8NwN2BinvBdHrDxHO51PRkIfWV+QeoqSEl9L5sk
U1bMnDf0kM2UDlsV9AJAzOKov9Vv3b2+rErDzG0pzU0LRud/X330fhaS6xgaXFfzFHoe00ZNiz35
6zA9VDXDM5WbhODe6vsEebwl2OERfDtxxUcYQUErDvyS7PoXF/icnelRJJfu5/qlWh+F8yPmQlIL
2kGr/VD0fDcGbexcgLKC7BukTy7sfiYAfWCI4ZDfGRrUYJo3pUiIsih/9e59kRXdvJ/xgisTolqW
YcSXtoRL4Hh3UgdZJoCzuqEcLjBVZDaEWn+4dCJNLKvWyTnMgo4CN91aabSh/37mN4WDMWd0uIvR
xbBTVfC06xHskXlM2IC25Z+eV2wQZhM+E7CpX+zhFBY5vYrM1acCXyniNrSKDGOUSe9Hj6ZDSdRl
3rvXVQLlGvdgShLryy6+p0tGan/ejzDzkoF6RwoDqp4qJqaAHZXUzqP/gU0jKNw6u6X9vAbwTs2K
0gQJ45LdPic2h2kgU4DCzcpqhCel9sAF9eMmjfB1/rzHcXt3bO9yjSag1nmHGvTZZlJBE4GMXD+A
XwEareOZLtqPmxL2RULiLomruu7ndEBwxapDFS5kz2Hqd9px+tf4Id4CeFL3hx0M8x6PcifOii1Y
WRqXD5HD2HCiTYr0ftHYqQd2tASw7d6MlUS5MfJocjrROpFYUWQkYFhfxB3rgRKLRc5OIGuQyl3Z
9icUjMSHcfc+xeL3BsMPPFGyG+vvVmKUhA/lnSgaGY5I1174QfVIv4ttOKuaJj4FdtiW42Vvih6/
qO2qs6s0ebVNIJnnMFWMaYhyEp6RHGgpozfQdS6DgDIixvB5o5v1lWQltIi4XyjtxUokqxy1YbqZ
CT9wmCNBly2hYSoKKPMS1so7kb5H8p4UdL3JXTHcEI6MujvHPCwFryIvceWI3TYMze1qruT/3bws
/qAdd78ZjuSDlsIe1jWjecj0AJTxY8MQiFQP2k9Dpg5bC5l9JNkUC8vLsFRI6OiV1FI6Nuq6jUTr
htCPUTSWNVf2ezehSKh3hOkHHT4B7lG7cmPtGN99MzxksjHGi6B8nVMEJo61DeudDp8KgggwV2ad
xk5QYSSWysJDlp1Ggk5UJEqr1hFZsEFGNRRCRRLTVY6v0mDEqVYzbxCPxRfMKbLrl36w7r1RCE2V
dGF2m4MTpLQP5oO0YXvp+CAVWIOp2aqZDwvZJhwXF8pzA7k5D9qyEgWyWeVMI31Yr0Ll+OrxiBjs
48H6555t7bDOFLXz9b4Qpy6ewt3L1+DPw5wqahMVrJMBm5dpiZMJbHLrtAK7qQDfVNfqUAbNqC5C
Ky2BDkxm6NKCvh5GKPmLb5RN53pKsF/VsVmdoia9UycVKoYpudsxIKg5JLRYXMGzrq1WWOgXywzW
qdU5JxAJYnAvt3vm2/0RMXSjinMD8oVtsj1HsQLMlkBPjB3N/1W+ytzpwy5LxdwEptBpJyYitB0a
KgxUaPEROK1LAaQCOXKiq8jH/nkqxR3X8jHJtawXSkV0dGoBrrqMuj04lDh1S2is12Qz0bdYz8Po
wAPc/FLXB7ro0xtWXIU+sv9hEfeWdPKl7stzHWfH9Na71yZK2ZSor0I47F3COfGTavqJtqNRwa5u
CD5pfRQ+4ld/cvJhgxO+J6mTY8ysTda0VjBwnPyzAcoMxrp//rRBKjcRR1QP/cU2HfOXlRiVfkgm
Kcamy9kVrY7gSNYJt/Dq5cWaiZ4IPgtMoGscsxxfXClc3VPdwidkI8LdEn0qHaKjI7AcimwptkSJ
66aeV2hAC6e9hT6/neb7P8IfssErsXkoifto7Wzyjq+Wvs/BjhwIrE0JW2XhOqAIF+lO7NUg2SDC
dXfcg/QKANpvqwDqzueBv5wT71l9zvMVnBgLHdBCAtv/RMy/3SBVnlXR+s0wHlPIlZIr0Fk8qPM1
Is9L+r3ZMSJMk/+MPsBdOqMv/HcHcByWHmhTEZ2eLKqjguNVQCciKk0a/UuZg//YQYSiGzn9LDGj
of6YNPRYl419uAftbL1K7riMA3eAF39grQuhLrokgCJxMSVQp/OxK+TYMBoq02bAf2CUnK4PzKwq
uAtXGEMF8Ipx8gZB/udG8XkoN3NMVUXYNvh406FUNQOi3mlgIJieHGMYv4KNxbq4HU1ZE31r9zQP
jnriSD5vcKKSxJ13QVI587RwYWYl9Jh5UcJDFjZzFssMNn1AjYihK6a4LKxJXJI8SS6FvR6IXwmB
OFy2TxNhUH8GOQHuIVEZpSFPVgRZn3mfVautXZzcINODgL/3poFOOD05S1v5YxvDxdRkVdCr6AAb
46P8FpTvMUXvmfL473od0dfRghxEXOQ2Rlwc8F6YBhpuKa+1qe3GVz76t6cKdNjYKadjGIKIktoo
cojf6I2aitrkbucXLDYUi7TGSMJTBmRWOekVNvJZKvwrvGKzOs6J2raxvpgzjTktbGpLDKJSq0i2
tZ0OJsU4LBgLa5vUZPcbyG3a7/l5hKnA8wGPLpy9oy8vCzg8TQgsfv955J/6m/NmjchFw4QbTJ3v
EZMn9glEqVQj6KGscJr2ZQybAz4+WLUl67VgrJMtPt6pJBp+yzwqioF+0s5ofFBfhTAUKLAU3SP2
4naToDmFPvvarjrWxRan9thdvgSRRLUyc6v98WZi07LZdyjsnZlE3LAg0eXrFSN3fwSGrRYDwtuX
D8LudqZPJKAfnhz75RLeDYD0PGbtMv++prCWTya+OaC9xWT6ynERaa5w7DsKSuGs8g+FemBqCrHs
jlVBeHB90Llu8gqk9z763UVvHTYt96rRfpHG/yH40u5XcmtsmSbKeyarlzHuvErhc+Vg04iIbc34
QZ1KQH58Ka/aLKnhBEZFPtf2x1/9TMjNXp2glRSnfPahvTMpc+fiO9L1W+gw/n2Q2dsirqW/Yg71
I7hd5u30S7nhttHvcUAz8IvvJOkDAmmplBAJRqZnOS190t92Ly0KnmraZip0q1i9PIMwxnD7tmEb
cu9HmqX8NIvBVPGoH+YpcuIJZDybvVc7z2+++7tgjM//dKkrBwvTfGNdzwjRiutaS/zDJvNzjziN
2jDjWZfb0zCDPQl1Nk9a+9bqvqSGiwj0XkaS+MRPqQHS3RIxGl6uVOn3OXREcDKdvVIMWpQDX+QE
l607bf0AkkwAM9nEZxjkTNJJdZLzApoEaGfz86nwKwQDj9o5PFG4cekULBsK1dPlcF+Pz5xvySwT
vZA8nVwTJlwOiT2msgJm+kPQb08ZgKCslQtpc7z/EOAhYzc4GGU33Wq0BtxdEb1IyR2Cw8cOoCUf
X7KvwGZKNxdST153m3QyQve28Rv0jU8MwwyrccNfjpdrL3KX8Qf+OTNyK0sJQ8lWmJlwWuxE/u4A
80N1/90If0IjhYENgLpU+AsKMnD4b3EKEkztbxx1Zyhrr7O7HNNElbwLkVYDuaK5zKfyQHZqz+MZ
0LMqjwd+dvdiCqroy2EWPSKr0DgKDijvEXEvS95FXDrRs5s9YHYCzWr1sSKEfsqiOvNznFl8aXsk
Jj/g0ZNAlBitDd4EsbBZMK4bdniX1CM/ufb7V9BkBU0Kj9xYH+iPZ3slR51PUoW/0FgNn5KQA1my
MU9pSHCeVdXB8ISs0O+Xy+Y8MRI4OJeB7l5iNv0n/3UkkmPoqx9Nprt65BrfiXdm3TlV4WBVCjvS
2UnLTsvmYMa5CH82nsC2AkSaqtZ3NwpayUrio/KgxJa8OPzRQuKrlT1CBRGC+rpkwfgM+OmRGxNN
xAy6awAH7CzPjypl8fFulrygdGrQSQSrRTWh4UYaA7E6shjyd+1+3mkKJld1fgt2uHHQ/LF2oEW/
gQPVG8QpObToUvTCHUytUK/SMplbd5xer5W1+40a9Bn2yINtaThAEnTNhzmIzKS0HqoBz3Anw3eM
zA6lwNvHskO5P4YNgrndjMSCzoG9mSLl8ET7wXSy1stJCzO2cwl36Q6S19fFWwLAORFx691wQiKk
xxwxovX2W8B5VcXWCKxFN4l1LRQfg8nUP5WkWPQSd9az6FcCUC51yK0VlEEBC1x6uQEnnxKtDV/K
SYuUo7KPOK7rHcdW+7pKgs57kN6I4SJkX6pzYjzB/JcPtOX6BdvYRSsHoFZVSqv20WsFfXurqhv3
uRpWO7+61d+xPV0+dRM//Y2Uz0d3se7EIxusoIW+QLpw8qHYXlJWD8xz9WXYzIq/uXkF1clmlHf9
RcrzySoHwgykRXhN9EJuUqvq38CxtPeWpEdgB7ip8K2DhrjPbilIzdRsxZt+0v7loCN3ZdvKqSBJ
XBysTE5lGM7xStzgfPUyzKev0Jli6DIxCBVB5wfb2muKCUqAmXPKYaL2rZXrEqp8xxwrGJZfjXX3
LEudi0oKnfRWGiY+Zo4BmiIBtD4uS8n7fJt6PSpcIuImtHUY7RPVQA6DH0F/HzteFFrNKQftC+d3
U+YOSQVFeoaovpvQSsrVW3LYyljlIostugV41OFrWUZ/VdvDoa4BabNbiizu9vg7yTJ3YJ0zqQSh
TjlimFznYYlZLEhmBen2GA7/rF+FqUOqwyHq4Q13EF9m6Pa7fJqUUAYX7wIOC0X2v8GYR+p1JTwz
q4VcKQdYsPe23WdHQr0+sv4ibFhPR7nrCdVhsF/mTBhIUe0fTvBcXZxlHdvQEhp25PxeFQV8d22c
DwQ3ZMmdezCqPhPDMRfLQTWtmSJKLkY8UKp9M30qc+eCdfOL5f8JSc2wGtH2J6k4N0Avdc+OcTb6
A1BCKz8qA7R2npro8gHvJuf4UQcdiZMyAfofKHOQWY5ZmCOvHG5pAyeCBLUCZAT5hQcVoiAnUpkU
UXKJZ0Cp/l05i//0azr97pET37ezBROJrLwK8TDcOtg134/j8XrKLF/XGSbxOO1T08hwPU3n1Cg4
XPJC22cStqz2ar2Eef+0gyhOcgtXYcCyMB23Hm/Csm5uxV//vlxbjBHRpar3D5UwwskBZ3XSOYwx
ZY3H1RPLhAj5fP+xb71ycNT965Ndbc+EsUmnbCFvPtBT1ALJmqMGCjjc8ghYperOFanfi4UVAKtU
MjMUKjFhBd2m2DKxbwaXWEsfcJzWtL6qVmukZ4OwVNT9xr6XpwhlkP+DSaZGFbwYQHaEle2QEB8m
mKXfZIZO/fYJs+bviB3blReCiNpn1qeL4aLxOD/bvg71fhd0yr++2l6dwTmmy/V9J4rsXa+VV4gB
LHEcMCPFajcnrfoQM9k5MJulAkCd2quMWQ2j7HXsRVKqUaHO7sj25V97a5bB0NN3L5b6sFAbvXpI
AOCxclOTstukplf1q8kQJUWSbYORc2nQNZ4E1CDN6Zv8wKckL+B1yIW6fGmL1UgDMRFPMG9B+JUP
oNEfai6h1yHyKzIXAjvXn6Mp820ZIK3mZi8kN5O10pKnLsvZWPGO+YllciM0HkoQ2CUwCEoT23MS
ila5W843cLqD5/8TW4OcQkvFySptK329Mr39/rhMC3oYfloCMP0Z3TIJ6DOW/SZg9arxep+6xBL3
IjkPjdipZV5NybR5VNlHDBo+6D+6legneGi/kv/A5vMxEMQuTB4X4IMm/ITw0lg+H3WCq97DDjI/
Ta0VnT5sKUQGW4rCZ7IiqQvC1V9Wn4G2DzsFZ73WvHgGQusCtkirY0xtd/UHzqidHQ4viPEyYlvP
cZsqx6MyvqRiZuuH9/59qcqiLPQYTw9vbVyIcS4gfM4ao/xMM6Gwyo4D4V8hGGoUKnb3SYUExcl5
idbWv56hfGI1MlJyK+vXdqV2vF0ZqirUgqpqZRHakCXxry2uL2cNVyEplvqWUuEXMJCwrvoTWOl0
2rRa/sNG4xFVJJxN6ddkWFZT64JqoLNISK+4b4qvy4/LDmhM9dSyb3umEi/JcmY2iyyOcJgZ/Jij
yzhEfkNgOobrN28s4qx5gWRETLSnaKdO6QORUdWG/Os7Bfq7UAnMVYMbSGF5Ns55lwus2uZvkRl5
G9X2s2yrYESSI+mtS3l3yj/a8cNDtWExn3E48ravCRB1rFR7zjIyRbt2uD2jYCbC4aME20DLfmCL
5iL6Nr7xXMyaL4lxTsnxwh2+N50nEo9GOHZ8bP35ILn0HByyCbWDPr69DtmmLL/yZTmQxUxzM5GH
aidqC3mxvu6MykFCR/DdY10Ss4xVzYAgBZYz7hMZedpkblgH/Srz3xWMPC2k5oEsKwbKC1jg+DXu
bu7LMWZZH2a9WqlB5+Z+Sp2wAKsrUdxlLSdnZmV7iCcN7Y/uLlat6NgLjV6g3B3pob30jLcKmiTW
xSoEFJqtnmk5LowG2er2Y8MclZ09p0EZEOTRW0dzjp88qLk4VVF2XuJw7KEtm1IM+tVl2AMfiteJ
USFQYPhubH3hJD7uqFH8Fftmibu/5VskSpmg242CEqudbLB4NCfkTztPTupnMq6cAOGbfxS4G4SM
zECs7me5QVAEXldWVuIwTcTUdBBhika+DsxWlNaH7cGLdody5+y6hmFmw56Jme7w+HbuWZlAG50g
enwnegScQ0IAJFq09kyss/I3zSFZmiNrQQ4FXAdMWjTR8XKYhGlB3huMXmAmRq6rrG3AY1WzpEgK
+M4DA5myAqwYzTeT8/YuOlt7BS50+bfcUEDYA+3oR7uay5d8qrbjYGyQlzCJlklYJ0lwu/RS0aFc
N9TPhaWxi4k1xtRjumWUJ0CdB5LHXmzBA6oQA2KIu414wGlPLfUWvjy//0WCzjeFHz3WBU2BFd7Q
NyacLWSRbbe2IKMwBzS6b8hQiVtOITs4kexJpUHUZyo+h73CawRQQHiCFS9x1LZ7x7Hzj3OQ4LZ+
GDAyKntwDfWKU9w2PBWW8phRM4NTCUs7dP0PpQ1X2J18y5kHKmpOIPGUse++fn/Vp0BwdYWGYbRr
6auenJh7l9jczUrOLR7Dd/ctq4+Qw9eIHo6hF7BwnOJ16lmzZEpbqe0BSDyh643qB5VkQoswMnrz
6K6nE5D3miFZ3omGVzCdlRwredq9BwODPpUAwBg2Stgr8JYHBQqaa4dIHWcTCORM/HF5Sao1L4uh
Z1czd0lveg0Li52wyzDg7ei+AoCe4FgQ0chkwgQlIVP1i6ZsQnNnecN7tNx4/FxXT82hVE7LNBmE
iMzHvSzjTPYbul9GIRgf6YB1kgWvBUCaBqwBlpTsVZ2EQd+YQ9eh9t5tTHg9326aiLYuquG7gOlV
SfBP9mYXuRAz5smZ/NdKYSm3kUkQFIzTVXDNoEN5bO9nD6lPySjm5rFo5CsupwF9ArzSHf5+CUzW
hp1XBqvgWsT4IkKJBDD5LAVwBqW7KNMjSWVhp4xZ8iPtrenyps05qwUuko3vNoFKpfih5ucmF3xt
RLscjGFYLO4VV4KJGYis73GVoiUDbYz4GPMB01iLXui/4gTceb6oQenbTd+FCFo+Uc2ZwxS9V1tv
ZuVEmFAWb+TmAqzM5YwQV1Yl+zMequW+ind9wwrV7GPiDAiqtCDZ7uoSIEG9+xS6a6/5bo/tsmiI
jx4yOldM6JtUhFqZoXgoJnzvimIcGn+W2mibADbi78Bm0Y2YxorlXWw2jRAgfj5Swp3FFRN05TNm
rJ3tljq1BbsiCFYrFbVRC3nHowrWPQjpNI1mXoZpL1SDnvIELEBYrVftoCWQPsg63HSCZKikrkOW
Q+SMW/jdy7jUkoA+yH1VugySTQUr8N2CKAROc45F8gqmI8+xzQbxiMmM252refmiQOVFUr15/3CH
Eh1Bya7Hh9kVvpWnwQzYAr2w3cQkXVLwdjTNQeLsrisMqzPZrIzKIfuMV+3YIjK0sh1si1lFWXVZ
XdWJ8g7CKfM5QbhjYyZfmkIAxs3LwB97kab0V3Nc+AB3b2WK4UJeWoKwon2NSg3lyauMM2LDUGho
zlcCoUi52CKkzCSdJXXe3yjml4XZOO3tHike4wgBA2X0i/bvO1jt74VXo8pvnvAQHfzcve7aSOH+
qNpUNQL8lGOqQc2YBVNd0muhYKlh7LjyVC8J08LoVyDCR6FqJGUswNJZidCIHuHSbMdSDwlJSO4F
hPKXb3Gd1Ij/qiLB4aSblQdg5kXsKq9S4D62Spu7spo/GI9Yit176GeHsL3sKWS+RcAGmxzS+jjj
6WcssKJtZ2CA0nI6buNgauJHfkbuj03MspkC/YoB41UW0dP4ytNyYPxVt+RAOV6btZaSoJuFyxSU
LrfKwpWz7TAkF3MFMVrolzKRlPtgltkDL6g6yHWDBPY42HQksmx3a/3g5BX8O3Fvaam+DNds6AXq
1ibNlKxasQ2GVhkUFpbSwtD56eeuuSLH0g2SNuneyD3RgEora/ROmpUkvmp1VYZbpi0P68TKkYAr
JMAVhM09hgH6sf9D1DoJzWH6mjiMz4fgN47g6yRLNuym1X+BLMgeE+X/3OaEphMgIFOabjxPyhsu
pYYTvqsaSDFXT6ItTZyzNcWU4g5nVmF9qOyBKY98qx3ChaQfJrtb7UdTPVJHM2W6dKKsDq4u0MMC
SPRKhFHTLqB2LDlXJoCA5xQiPTWW3wUN6WRboA/sBHJntxHtxQajzuKdKwdiIjf2toUMKNL5ArSX
2XyWHsrjRemsJUzP16NtoLE98ux0TEqi3OCQ0b3NkeMZvDlOu47wtckZXADtLdeozVLXZm5kJuVT
yeztCo22nnYuuYBIYEcH4r0Q3OeVzZ5k5bN1PtWdM1OC153bb7ZIKlHIZlNJOukFh6owHip8hiGE
AvLkJn9oHngKPuNLXpWF1iwXbknsAp5YccpLIxz+aDi9sZYM0Xi36mVitjer5aEkN6qaqcG2vMuS
xbzBrID6ORLOI3GkzKjNk7AbX/+jxstCoAf0c4avKGVM8dSlsSs+6V3THq+iyqs8kYfe8LmDR0gV
bH39fjoj+UUPdycwQpP3ecOV7Qp6/l9XeVnFZzS5vck6a1tIHAc6QgffQIp320y/nlCv0towtlie
mw3/fexwVw9+2SwAtJBml0wShDhut0kbj9hIL1XbObOy2dk97d4EK6LQDFsAN0QI0CHegcVxwZpu
x2XxMg5mk/zVW7ZFD+6TEuJrhN+Fva6B/tNZD3KZrZM595Ab/MzcZx2fox/7ayAsrfgeNIqjy2B3
3K4Kt6pgKx2jNOnkSbmuYloCI3VjYlUgZgIdTjynsxOAltRI9zQNV1X3ErByPWRiGBmEg2P4HuF1
zxByoh0MCcjR12HuOb/QtiZriQrZM/nZ6ymyxJSSDHgWOJADi9T5L5H2n8KAAP7YRYIqT4iu2pda
9qm2+/TXcI70DNvD1QgKHDS078YA5hzJW2mveSRGopzgK5TPaTFOSo/4mZq8Hh2SImkE8TehYVIs
ftcOjQpttGvvvsekc8xt9hAtVIVPK+IszAwfeDbPfHhRU7LHsA6b2N1sIVgy/1WiG2w3CGKsDzz1
7xm7s0TU63LNe1ndvDbHsdpKGeL8o9EWUvkPQ5ptdmisg4HB2wB1zOStAnrkSlS5+Helq+joOdPa
gzpk1G5kkHnA2ljPzcCby+a+T74EJpes/82sS6N5EKmMsmiW4qPhCFPRVnqZEKcvAlqPXfaKrHvS
gGYjq3hLPGe+G848ggc/DdSf9P3EmfBil3zjh/XePUEpRyply0mJ02A7A8GBI0HMbcWY0eFw50mD
TjYEkY/wOkAB0uWjuT/31UEb0yKGcFKJvjpBDtE22RJ0fToaWY2Xc7nT3R1rYMVeIW9BaS6EO7St
PAgGAgJApLRsexJgw+BjNkenVIg9AzZE7HEV2y/XdwZHzB4O6U4PXQGJ8+BFlPgtaqgoaSdnb4ez
uSFpgvaRrpM83BhFRqBwCMbfITnEj49TtjeoTHqfy4SwxZ7TOaITlWfcvbqdI0/2FTrPGcTLWpcZ
/GiGvtoOpNHK0tEZ2g72MS87VWPaEAaPGpNsLM0eKmqBoliWFmfKQbTqG2+t2XqQFfJkDjJ+Ap8K
VrPK0oWygxhVfv1orIFtBItt+jbaX3yGgASy+Y9OnlFRJgW76ajFcpM1rv6nvZ6bHO9J2rny5dTz
hJu30XP2lmdVOOzvti2IaGWd+TQNP4I6Ovwo+9TfU6oP+GlAtx1rNs0EQG3gpzMMx6XFTeYdbPZS
SGUw90iux2p7hvC3l96UiBYv3TeONmFhj3zKM3ubbC7qkzdnzQrD1Np/rmmLn8qqnT1pL9bfHVzG
WDMu0lCOFOoL2GDdfS5j+ewBB24T6hCaMzpu8yjlx1ccuB2WtD26+jxP7wadnHnkJ0Ra02Lyqbe2
fe/ezvNQCIvy3ze+5itlEKS4EcrAdGDToD3JgFpz4trUbBmS3gJBThj4bU3rs0icacmkMIOMDd0A
BhjYkHGra+yDpC1STy0wp8HJVF7ccy4N3rCW7fy5cK9mt59JxYh3Qy8MlQTd25k0oKiREO19uIqC
nzsNJwY2YNGa+wg+MhDNQYbB4zlRymzB9PLnNW5sU4htku2DFHKLwFknQlfRaiashOcFP8LajSDb
Qw53ss7qlgQh26T7tg6kaaTg8DmQheppwbWsfMo5boOkDEIHLHJMPAfwIrP9V//kO2naH4t5V/Zo
85QYaragDqvtvsKDHjWUx3mTdkxYhwguXKVxgKYOQMMQosA0H22X+Cvx0sgLVi5BoTkCTL1+eVLS
RWFDDNaq8V1U6Nc5s+t8P9xlqg6vpd6iKxCi8X1Q+q4mzGkp9/LiuBYFMLPtb8y+ah7MkxlmdDvF
97EvuAbPjsQHJcfmjvXCIJDPmgpju0KIqKlaYThE0rQeV1bWmCBQ6G2uG71T9D5Nadj/KfdARBP/
kFV4yMXdVi/C7zntr4rBOuJLpXjf5/LvCXBc6G69XHLD73ZF4CZV3p77d3eLOn2Xjlv8h38rDYq1
x4AJxveIE+xXuP7mYHoUOXnPYsz66aToSyDzLj+PH9DHS914OumsAELoqcvMsHA55eFQNkea+YJ2
VOycMcCrbXtbjD4mWKMD9SCxMi2Jww0TzzcFuQtCdHC51T8DQherRGTVU6eLp00VSteYyddA/fnG
WbBX2LBx64jzEFbxJ+/qfq4VnIcqnFiJQYft7BzEIhVvQ9elD3SyI0xJyjptlNa+gb6SW/qCGJe8
3FwM8iS4mQ5/zSRL9wy38XcxX4eMlpXsAbOzpZEGrYuxDwd36jQnduINkR2iFhMdsJmopmU/oWUJ
lKPOTqHaU6apvOgDf5nZsYP6fu649LsHyZtfNcOVQWh7KfzTX53vPLz0Hni4fiQg1CFmhW1QjjCj
pSjcW2y5y3t25yQao+3PCBwU42n/vhgfzpTx3xsxaVndMI+WYnM5yAg9pRZQ0u70xsx71fv3Fzci
FH3XHGDuxTwwN55a0CA8YMlmFzZUbwk9aQJH7KHzkfEktKbxbe83HXjWk4fwoxbJzJEb4wLG+vz4
zW5ueety4e+EM3kYA2gTY8rB1wT5hqxncdxVrSdcmEL54Z6R2Rc3rf5clKA7Ks1dpYLAXXA278j+
KwOC2RNP7jws/Zx+plKxDX3ffRD5GJoZGx7ARDbMB11LXv2lVjN6z5fqjzp4pDz9gGIxK/fkmYS0
gJsgivzQVoHKjBTQYTK1ukki43LGQXixwyqVb9no+uujQ3xqKBqrv2DxEEPLb2q2kxYvZWklQgLT
0dhN8IXZgYz/RMUo1k1famhoesbYPnQNEpLmhFej1wleVhxz3zh6b8tRhHFkTwSrxMr/9a0S0kOF
/3DKXn3OGaGP/ykZLKA59wwerAwfLudu1VJ7FTGwch5H2qN1x58CQgOxp3/ibPVJm7N94WwnLG4I
iRzoFCibqZnCLxjgxRQg+KVAV6lwb9OZbx5v7BShoeAoOH4AjJ49EAKyDQzgWq+FAh4xBFL23z2p
MAxmy0ebz+EOotfl6s5BCGYbT2ZY5qU+rxX1/u3XPhd+BfzBSzFbnjxogFMv52W5wMAY+bu+DQGq
JQokB+dcAfR1PysNHcafFlWrhFsgVzkX845lo+j4JLsEk5IKkWj3xzBKJScOvFipFsalf6QR26HZ
Oy/sh5WQ2PEFkmhkoxBzmZVUljkQwgtDOHzSG/qvOTti0wm3nxWDEcJg7E1Sonx1BTwDvhUgSMMm
5R2VqEqPd886YaFePofz3gSCesjF3/6Zp15rbLHLb0cy1AKBpMDOtOCBapaxBG26mOoUYoxL4S32
sgdYKPV2XcnH03JOqrANtAneAoBM9xE2CY0PpVpCxFaHeRW5pz5E3BKOM8R1cBnCS+ZL4yICruAV
aXGQh5DPFgj6ZoOJpN7SbQzfxNITm69h31EDPrYBiNfdHz4z1SG/QqJuZ/tI3pKpibzsS2rmdD7v
Iqz+8mDexjzuEOw0zUq26+IQ5eI7W2KNMrnTh5sYKLp/wpv3fTHxzR1DPZ9x2LVNvXpWx3C8eJ/m
BkqIbN55vtYkhCNqxmWopWrx2/CcfIZ2es2Dv1YEUZQthLqKM2JiQr50+/AU/SbZ8HGJXkJOtkJF
u603kHnYFWIVC6FB/bSXiLWafn9raFdqyjzFz6oz31kwMqfOxGJYD57YsdAJsEVRRLIqtUbaFk7e
2p4P5a67BAahg1c0W1ewAT0sP0dZL/7Dk+VBzkNFzQcz6f1E2N/Tu/0EbmJROgjp8Mh6GaOyjU2M
cPRJRjk3IDVyFz6lmS6PLQRHukHKtHJOuT/k/mGtoc/6nvTZ75/MNm0brXYB0TO7Q1YpcBpmpDLh
D/BVL1w7nAa1wmh52axZmyUNcpW8y2LUq3dGtQZjPpLEqTHLBHMlJxFX/4hMJs2ystYCT/Glw4Tl
nyrA8GcUCnmO+CP7Ey4rvmzmX5RcI4srUlbAFMBn1f+IXaw3tcfsUJeeuWkSFoZdY5wXXlJj73aj
nqB0BLCusAo8rSeg5VfJDH+ao9Y5CSdVE9lHqto1vAMoPxwXtO/M76Qgsk4MFeEPF7+gjEJHCOm8
b9V9+xhrbaVYKQuoa1F/yICvTI0GT6/d7Hk7msmeQ/HEVh9BhhHbTG0m+XMagO4oGEZmTzmui73N
eSZSHp38uLPQxr2JXhBXNw1Ua3jsLqEWcRuqogs37OtTPGFNUknyVWrKFh5isdnLQPo5lzaHvOAz
CdXBCCQUd6svb9Ut/hHyByqXfLjxoYTgalQdcDdiibxNdfwWWPlbhilnsmbNGVFz1T+THHJkHsHw
U0vd8QtxsHnQ5fEcVVhgOR6Tioxo2RBIlttU42Xuj52O1Crl+FYKSvCxBv/CXyYVJwznmD1pfB+u
NmBNIdtsOocnU1Q8cyzhrmqlXkl2gp11YPHPFg0bFIvPGMp/eSDMTsBytFGv5XzNYJpNUgrCInIQ
5lOTuAahQOs16CyM83qkQYe0/3OFEWCsYM87EKJ7RLI5vVM3QRaYYwLxmwkh7yGGSWBplQLjxrUe
3KsR/TPrTaVOe8uipxG5LlCMhP+sFFhPOqyz5uCa4+Ku+vbhDk1ihnE4khBT38CeKK+sI9rHySCB
fQMShJA2VYBKuxUy6+8EwdgWAVKtuOtXhmexn4zW1b3WueQ4WiFHKc1G2G7AtZMonEmeNEz8mJ4p
KlJBVY9qrUJs+ILj09uWcu1H5TtzeEw3Pt1fR7YMEU/J2cnpEWCDOfheGWn/npWeF4G3VrLZCkIg
I4P4CNliTQ880YT2OQ6T+5l4abhAOyrspB1qG77MCBfJ1J42+kmLehjyVx0+u0n8IZ4Ul7bwSQAq
3OhcZPHTl/eJssj5Iq8QJGoFVyDn9zN7pz9u+SkdLHYi450WbHeopKkaxZ7+QQOwx8gnqvnziWMa
bMFz2TQ0gHDtHi9S91IQxKIlpsKyO+z1KmTbo2xr/Jv3VjMtXBzdWVClhXhZYv4Ge+w9DRX05Rqv
uKdclDza7TAHGy2jf6mcQ6fIoQ/9lauZHMozanR3VY6aAWqGcChV21DvgJWP+JxRPbZzx5B4Mn8q
6FDr51M/Abx+JEekCfdIVf18alROvkyimL7dMLAQPp76lts8visq+xYJYg4G97zV4W2KtfLCb4LQ
R+ctcoCUApvrfN6EnbLUCifCPCD5lV9728ms99XENfwehJ0FmTGTl65jgbclJzKCu1sCElFZceNn
iSrH83J24Jr/3qI4K4ZF7mkEyRCTTrpZcy/mbgXPe00x1bCE44RL5rHlY+Ng9dT+bg0fjj4yyVjw
ycjVzhgoX5TOHFL6VQGCtb/NeSjx6f5vBYqfcW22QXpN8QG0+7n17UCQ5+QHdc08kqRLtBiy+hqd
AbUiUAzhVwrkXzEegV/wWZhRfgSKN3RBKNBX7ft8mhCypYhI+DV/Lrf6EEv//IXr6L1FqnWKwmzr
WvaebrJ7tSfKi0TVk53hG9e4VYQmPEW6STaIn3HsE/1DaDDx9RGCt2Y3LBpjKPYlQ4f1GzT4A1HA
dJ0cSgnHcYd1K1ecciUQe4JLYo6P3MchVCCmrMHI8Y3oXVQde8UfrzzWQeL1kdexSpw3A8fQcaRw
6cKSjHxV9bhOxz3ZCPm1CUybR/ynziaLLM8xHIiselOeXeqeN+oT/vSOz8f1rqGnlAXvzPrLk+Nv
XptWxsWaXP4/tNvCwJMfh13XRt+yIQod6XpF+oUpGNueJR1LeN+/TNbyF7KOzPl9KySrhuUf03lS
fHzVTganePw+ccW8dJ2wd4x+pHxQH9aslo+dfJcw89Qy6+tmhEP1lMjlJ0Cvs+Tx7jrtIhFtpOsV
0YChY6dBfWu0hZcZ0XuGmCbYZRv1MbWbekaJgkwQ+4Cz7MU3nl510mFthvn4iwMoBhy1CIykiSn9
4huc/ZAQ6zpxDJbtR56/WXB7A8E7CbeHDDl+Bz/oDmNt/y1uGLrhVDq+X56NoNXtky06SlsNiNLT
tQrSCvDSWHw6Uh1gEgJpnGUxcNzB6bBzwg+RcyVjpQI7JMl1kehPjAo+lciXh/WbiVaXqa9D/hjY
v3QvjMwbK8IMkIsQHesDagHtL3oDF2JrBA1g6L+OeyYOuhoqqUMHjhcg5Oa8buW6tOAkTFxqt+wq
VxuQ+rSdIdk8RdtahGwkwtVuKrzvl8Cz7xhTnrqeXb88Tfd67PMBgatu7N+ABZwQ9/kIAH/12bfG
tmTVwyVXBwKjGXXbAhClH85RZ0wXbd9ErDO3H8EqxCtyUyh88Pw+wW0JmBCvaVXKnH4xWqkbPOjB
QGTgsLS9xw8HDydYDozUYNenFIaNduWTSZ+svQbuEA1Z5zmiWLzFdvw949WvjuGStoKV/N9bOtkR
AgqtKVTT+GyPOOJ1/s1ZIVPrPzrp/UebP6KvPC1uozfVZe5uCQo29ENXiyJjuQZ08w5InhuGTfUB
D65lY7sW+EHZz3X/3ulrmSwx0ggPzTncdgWR7x4snhIgNpD3+cjeKggudgkcl4peGKnOHcicJNC2
yEyoAISLx+d7ZnpEKoIMgDfZlzivbY1PYWLqI5oZ+n9cF/NFMIYbESwPInEhgBDwphqPSaHKvNw8
TsMkGUWKxOGfb46F6Lax1kikeYfA8Ip4DgMgUr9tXLJ1OrGY1MRSGtKeR1Pqo5EN5TMMlIB/ctxe
Aa65Lb0akXwx0EU/arTq78JPlFvQzXLhpTQpZhm+mDMwgmd1qwTOKJNi69WHDCJbIPhpkfbg2dK0
9EqL6hfZtYA8j61fSxdtcMX9VYFun1bJDaKR07c2pPYjH0EtdkvutQJafJsbmOFQ1BlBRRtibm1X
851EKMlGESd1073GpMzkr+tahSz/wY0pteP/LbytKk7QWImqlVbAqhLEIhO0ceIg7qoGwMy3iDJ3
RInYql1Bdx4hDWx++u3OUsIy189BeRRrVYoj08uCkaO3Jm2ggA7/Kk4IZXpUllAS9bSSnDxx4fRS
PAtNARVrLDPm3tsu2yjJjYZwt+1UHjV01jdWwOPI7MZB3t3iSHb3E9B+GvJktD34cK5kAvB1BXbu
IcoYGuW5Zr0j4/lwZ4XEM1rjMcPMIEOI066gNcOPSkVBdVgCk5Vo9i/314pXU/cRAL0BaHAa2LrJ
eklL1ZYb8Iie001Q2qwJAitMwRyLKvsJul8kjDi38sV8b8CWHQiBU6yneZzM9VPYHEkDz5Xz1hpz
9wQQ3xAtcrjrOYLzFZIRb+m45c1n+wMeL55cBRUbWo+lKiSlaYYWcl1wW+VGgtdyg9pouLud85DS
J+EwHflHhOzV/w0RWHDW4N73Od5Ed6YyIqVNPid8CwAYZSm6mxDNpb6ZgMVTlxHyHKulg1XQ3f4O
J6FCbfpAplBs1Ai8ypH4ZcdMx4plMeChnIq0VTUQWSuRpwP8MsZE0CyvXJjM2T2Mfzb/pC5T5v4i
byg5ogMmE13nE9iTvEc/AadpXOV1w7HAaV9uup47i+R3xyzqa3GdWZHAgHw4OjcYrtD2vP/cJKym
PV4m3+4bZmMPkte6X1EYbejhnK1pBs50TvHTO/PUUuOmx6WiT3EOs/ly7QvAGnfd86ZgHvKNqj/L
RpBBDFM8VoxEsorErQ7w2ZZEmXNklqVcAYXK+CvNUBgKj1m2MtZD9aox+BXRKbd/JdDeYOosujxS
lbGcNa9k42WCvpt7IXhqN5eA/Zvi2T0TSDHyJJvfXdNts1YU2HTn8lFUjwnOHhfalH/B0WTax19G
P2tyqU4VTDHHEIJ16X0+ZDEouPe409TxOdAKi8deXE2EZWEl+mTfKaQ1mXSSf89Z33jwAA7KmgUs
2CxM22K9bB4JZb3L4Dx31IwrjX1uQ/cHmfb22qbBAvCA/zDLkUQMrI9o4MWTKVLCDCFtU3kH/Zye
F051NEN9heLWi06qSguLkttdZ9S5g0prW6maeKtVJBR0MWEoY57BkIQ/VkxO6SHNhWDjo4o+I2px
ly4Gfpqe9KyArOi7XMJHYyRm6RRM0+DZ4Y+S2K4ZTj7OL2oTBUgHhgW8Ng86Rgsh6dEWSDLLyDF0
g6AeeS/V/gXd5wqKPApmCEGIwD+N2vXJLqrVIMOssDa8tgwLR7rJLcOvy3L3Eq8HWDrn2ZD8O63x
Li/7jSRKKhxzCOY5wDrYIwlcHnvgXMp4EzZVBi4wg74+7Qpj6sbmx4LGFHB7MLON09TCTkGXy+LC
Dtswom/ECKvYWbnJISmxe5T4goB1jZR8bIFJWUtGxbdukoS5o4axu5jHr6vjC51FjmJ/62QIThG4
SqkO1+k9zwDV7MsDTVWEDDRjBiltRvE48PASMp7KcIRfifhcbgXtR0AKHa/Ns7IcXtqNtLspigoR
eQCsv8ZBZafSA35huel7lIbX4x9rnDapCf7GXrJr+s8Cme4U6oHzwO/HcF4UwuzC7pjDjsCoz5oX
Byinm7jW5LJ0VibcuaO1URlN5v0iqfPM4Yc6KsiU2/+/8s0o1LhfAXkXN89SPQrFwizcbdePUjYu
yPwXklvM042Ufuz5by0yYHwmvL6ni7nSPKaJSJrSeyC5AusjZB25Lyvm6YsIkZBe8QgR6gK22u9E
5+qXYXdnCLVAhX2m8PlDFb2K5DeoUbVWphY/j0Eu8lgtcceQKgKClXkjsbUT3QL7G5nNkIyGj7L4
0tisK8Fl0C2u6DsfCG9blszPTda6qeiMAPMLTYapLgvdbtl9tAkrH1VmNN0w3IUVH+uHlNJFnTyq
H95r354kDSb7yyhV/KnD8lcw8YOq0NK4I2qo8wxWRTXPwFdJoOMxYbCIFpMJXyBEkTUzcTtNb/yb
saLx/a4A1PtAJUUSpPzQN1goiS3tpPXUSnjUGVHKFg+2fNfC1uvncf9ISQMIpjN2CEVGEvr5Fm8z
STeXqKjvHKygDCrDGvTQLLnzF8OT1/d6z7Cz1TcOQmuBrb1x/tNOwaJ6bAtOmDmVmw9nFtt39xUM
vtFPKoNogzo01SgoSSW7Z/rRxAuBBaGZK6tYRO0vbDGeFLIM6AR1J9N9a4a0jjk8heNHBOPMR0mm
mhXuO7jiKMy+4hpUh4z6pJeKYWOAA+SeGg84QZ/VV5sMHZWIkK9hKm5Qz9O2RrQ5CPxMLD5EvRlV
/ayBk89M2zH7Re/U60zTI1fpdpxFPYJd03oz24xFAhe2vGGjKU7sr6qgl0EUALd7rgw5XSrmI1za
7WkwmejQv0zGGgm2dz8QxABJCIh3rCfmOrmsGf4Do3mb4JUo9mRvFmLJIlEMGRQwMb+57NdozP2u
4fEFODUeIAdlq7qxQIRTjRQ71a5XaFH++BiVhJeCUceVnkp4X5XfIeMd/F4uiKJWlUQXy/hR1fgv
T7QRAgGPsuV/egp78H01wcuLOw0+QVdsSuRhCKubpW9fuSIJ/DV2lFgIrur9dcTrd7dCkZUEcIht
TtSJUIqU1WZJe3dfHFug30ydgSxpc5xP6tZH2OuwmnR6y8zpJIEfQAFiThpbqn/FhGK2dF4asWt1
nr/SpZOrfQaiSwbHbyARIGXAC35pLg23EdJp/MnJMeGmBHFOkK/WelYSunZBEdYKlr4Eyyv80XSw
Inz9EQ13z1u8E91lU6Gtfuzb8ohx+o/kBKRi95S7nmbXVF8RoTb523TTAPqlyoOtIrPLhGNydebl
v08RTIoAazJYldW2iHTgUMDp45eIywAOOR7259JOUSL38OE0GHDZfo8NRwmYJ0X9OCyQp5yX5xwZ
CpuqJo9YWqapvyLWVP0fM1JLGekzPEPfqSp8RzP6jdaxVBqHRZS60pmnVfuTwg+L15hcoJyvvMrA
JWx0DCjLytEPQQJ2zZsXx/ijX5zfOpmiwVxKSwtCbmVAEkCB0jP1LsCilivMpfch+YDx8lTZDClc
EWUVKxIymzNaC7UXInqCp5Sf43IRxnVESGdSWLQ9Ey84yeYBUEnOAneK4KCNcFFSRNTDwGffGADI
I87qh1uQfAedvAXA2jP9IKU6tEuTw2KEJ3bIWQfFRd4cTbWIiavzkZGXXqDFYL/4Zje+FRsTmvr7
PEmdPzbHFv+hkQavzrM4slDFHAS58/ZrJ0+CC3+obOzxD/jAduSeLfuCXwxWgRjr2fdEI0W++Ls+
/TBfxxNHLLt00at8CMcPkm6x9l0q4LHUxZSYAcVszo9vU1XSuubVzCBXV8M+Unm/xZNhUhUWkZMJ
ak/so5YvEXf2s28OahQjCSIrzkBFVQWw1qoIZAySI7wvaMcwUXEMwQcM7yq4rnC/CAYh5oaOkb0j
JGr7skLsFjOE3qF9eK0mvT2HAyUsIU5Q004qJCBnbBdXGrKJbaYyGhI3r4C+2VqqlUEbDnN/nR96
Xol/qTyFGEE0CrYrKHa9c6scTpMHhciI5I3biTbN55xtH3dVNdg2t7/7ISB6upy+2pRZFl3uwMra
abNp92paBZP2tZwDaki27TS/ckRtIR5JTpqRnxxUfZLHkwoPsoAuqM1BiM5qdCsqC5gaVSbf3Yj9
sXzAFFo1sotwJ/ErKIEULQcPmZgTbQu36Stt72sI5YiF7b/oemU7LeUumu/nZOQulMrYMH2FE5dB
MfcAyG9VqQM0wqFrLcr6RfQX59jBI9+/k0vOd0oNmiP3i0OXPVUsVnrFm9hdRtP5ql2Ght3G3W4B
fOpKQxOCA22Ki2mun3dOioRtwdLgxyVyGk8thAis09An101BdfUnxMM/trf+L03KLeUMiuwW/LMn
9qRXcHyJnD6jIEBggNu3CnaYw5GeZdxRBgcON1Iz36beUk/LCR/cWug1M6Tv9dOldy/06SV9UN/Z
hLpjnGZb1CvnxwLenrH/Wm4PdF+Z9CrdUlf4vqU+ONaxOthhP2algIWl57OIP5ZEY/hc1C6zV9wZ
+tJEX2L6WhsuwCJn+tGWU0UZIbBojz4jNLVNMmYZJ6utfrOmhF0g8Ea8fi8BD+23LXKIMU6rtFnV
02Gpkfebd4U24Z2ytLA5KBJtslNLlZ3xp0Rj85PwruwzfS5mTdpYFJiUkYrIqdXq6n9eag2VzmFA
v8yqXPbOfaMxomB2cIDfsoUtCFBjecaxKmLj+m4nDx1W5NSTUMQ2FpPtpkMVUSUyx0lDlgGRWI/8
a5JYkNReL7L4vsjQ809B54x92jQp3SYpiZqxVu4cOsnMZZuE5OKAA6vrKieViHDWJ8OghSE8Z3dq
h7WkatBfSMTsin1uZ6k4T7F9HWS56sk8N1kynYetxix+JU+bnXixMfgK6WkMsfoX9NepYyJ9uxux
gxtklP/Kis1aaXcVCuFOpOCcHyJjLGJX4lT9pnhAKyooHg6b0byt082Za79AnMg20H+uU7czPglj
epcB2T8lq0CSRtZHllNTzCS+csGtIYu3HMCP6FJzv29JLONTt/SUll9jJLhBi35R/+v2Bxa9f4k4
r2LFI6vUuFTPy+NYoM5mnJkluKdkFmD+s+4tHm97QqAemgxWlWApP2VQYkrb+a+lW9x4Uqw1zaHf
f5x67gWiMVrPBYZChf4ZuZBXuD9Z2McrVRISIxh8s1IoZQigGSWh+PeuS1TYy9VBDjRM51htdp62
YegbfpDtINfNThSqogJ9u1OETzX9pL4q1x4PeKnC9Fz9ecAy/aehtLCnCnsbk93IiTJT5JiA+/K3
3xTt/PxKPFHQWnRZedLeQNrdt90PU9/og9mITpCBvCl7duOzH30/qWXDWjKlNN8zsR6AKh8we0Gk
/B/ku3UKrzg/MsY1YtYkSfl/hhI/ZwsubdXpPqXgQ+PsH2CDLlHyWJ2YMVHIeo4jI/ePgOnBw89X
F2Z6JCX+1IIp+KcDMrMYwWrdKG+i3aPvGGbQJac2lLD7KsVzYt67MmQngVf/E5chizQzuh2v8MbV
vmBmJUE5fgtVokvnXLexPK3HD1XTrp0YxSOhxrWrPdQik8p7w3qEM+REd4t9XZjTnUGilys/IxeE
EyF81yJZxe29V3RpndSwZESdsA1VKAM1/BQZ9JKV++minVKso2JwZzmMRJLtfZWUBOjGRFC8OHLi
kJ0Vi8f2M7spZpZLDefKhUqcZd9YxpXsVmbfQ3FKb8rhIgfuTWFAok1pEMatuP39jURuQpxZ8MUq
LDzS7JOgpG6VqAOcsM9N6bufQzCY8taZMA7yaRqa/S8btVNHet6Ux/8pOBVE5GrNc/DreFWQHMRc
ToWF05/r5P7iNfJPYrEFTPTWdaMYtTUkVKSSH1iDejc62oYhivhl6QSHv/03pODzRufHb+0NGg1J
OjL9GDMssNu/XoossYiQTVGKFPe5H3J88HPxpG+pfuq77aCpaqKgST3D4CQyrV6ijJ7rSb0iSeAt
SHPPuvoKtR4spiAl1QKJEwfZ5aZD3p5312TsA61Tfu8Art10lkX2gk7/SpyL+ku5DSl0MNEAmmyZ
LroNXyHiY8Bg+EBDU268xVjjZZBXcYDS19JlpwSp1OcyCfRpEs6Pbwt+aGJVH+5k03j58ufx+RB2
cLAtZbqHnbQy7FzVCozrRudmprlKnrE1WZBjxUEa7IXjz0U2xryDoOCrLm6/YYTRId8MH2Z0Keiw
MTJ8OjkQnNtDQtl0Fc7aGmH4MpL4UIGcnAI5DAHF7K7o3rn7bz5REifucU7vWSuNGWcJK0LajRJy
kAmaHz8uXuMyZiza8sC70PFJR/pvsyjKBhh5YiVdjBT0NY4JkeFMGTCTNdWrae6brNiMihMIS83B
WcZfOVH361wZ/BXJq029MSCUuiE1VuwkzxQNDKtzipzEpQD4G9kEo5NEd6RWwGyzyzeszle2UZtZ
JD5NFGTxUax7tYFoS9CeSk+raJFrYXgsBHowQa1+A25h7S12JR5ouS+1nlyiLQwuwFwB0wfhoP4e
u0envjf0nYqriBrzYC5QagffcQZad0DZWxYPb9pc7ZcEQ1EN9Q13DrDGEe6l4UIcqWG94tRlW/J0
ZLZJiwpIG2GRUzETEFX06DBAniHXuJ8GkIE3e/2H0PDeT81Gspb2+5wNrxBhhhchjHalCLg3dSEA
ckIQuOWFDv2gqGVpVshyZGqOsn+u0BtwzRyB34nZp6yeXBbHTTcJT2g0E40m2z6+4QnMMcShQfxT
5qVD0B1hUagLhGG6r9TdLmZTzPGxZmTW5VW6RDhGEcSmd6XsjwcQgSXTy/03j+Bf3tpmDFPVfR6r
mnsUUsupR83k02Mk3Nj0xaL/HfM/TaXW0uBItDxZT1c0pWy7O7HLvO9wF/QcCi+sKENDD91AIsu/
v5ML/DZrNGX3pqYGg8QOba+/eCajRsI6qKn8BPgcHed7YfCHRAUoGi2UrDEjOQPuFb/xmhVcjtU8
fIUr0eQCoMvuuJ/ctRrHJagaO7VXTJV/EzSnvG4qllzhdDYrAPZDaexepjd/xoiQ2e3Y/AFwonvl
Zx9EJ9WhELAx0CxoNVKe0JfSQF/xy1Ve14hFEHzNcCBonBBx3mol4x0SidcZttWoBnUPlQZ8+FlN
y7fp4osqsg2wd8T+IJxAgR6G/QhxTjbuVJdQBZi1w8/5evzVWpB0rPW46JjsNpNwmALjqvd0d2kR
30RHcLWF2oSqVhBhycq62MOtl/UemihHXsdp4f8W3mBTjWNa57NhvkgA+sju7u2ywG0FMdLXX+eX
RzZ5lhhLe4g8RX+YTi9lDEfUBJ1n/dhAJnbjTpZ+Y+E7oPqdruBXh5eN03fuH2eSEUI8PLb/XR/A
zuQWhtB4CyMjBcZAMS+3Awb/aH8bsC6yPOI+CHBZ9o4PmA2Gmflt4CH4qcJmLGyyjp35S89av03C
QazFK4xUstBhjyFffednwoN3QDXZXlew8wskfUB96Qb7wEbGoNixxQVSNm5PijbaHIXSOevwvK2Y
morKLIkA704BsRyGX5OuwFnbIJ7o4JPM/KdJAFhWvG5qrDYc+/scI7RxOvzboxiaFKs8wbM61QjA
6hDu80CRB0c3KBJaPFDLcCigSs396iO+vzSi6ByHi5zivx0VkyRwDySyZImtmafAkqxmkuE82Fzo
IbcMCoDD8Js/C5S1xj/COiRDj8vUuKHDj4fEUQWHnpnAKVcNc/kv7WzJJ+auqFvxOf03uqnLPAHl
PrTMe9ebe/Klv4bGgXfe1aFvOhC/7xjH6sQOCmPiN5NX6+DtljEFc0rWERjH6Gkv2HeAC8d8E5hq
L0ZzYrFbDaF0bJslIThgNbT9ryvY4L8PlLCt80PBnZd0WDwEtrgGAdsf2xI1YeCQ3DEFLmwV0J+o
R9o2Yo8QqZtvtTDs6Z+UtQoF9DDygp+4u+9t8JNP66cF5zvGVKFkNK/zipBsL5scMoG2lPDNEG0I
gH3mFBmx6JJ2rIYfSI6nfneSWZpidHp9PF5cC7P4Q9SrWp9l/abNXptyvfP16EJ++N5qy0y8zVqV
0UXXf1P26iCS+GrFyN273wy3POGitSYWvSuulRh1nhyNiKJ0b8I2u4ipYvwyX4OJaZBUqUCrx/Oq
8haAwTmM976pWirO+nh5cVxEy4RDaf65ENz8ykTMTEyj+oTGefwCNwk0ayHMTIXZOHqmC3Q7bHd3
wE3NQ9Wrqegyz8RLrPJ/Oi1VhjiolHQg6lH0TpGcaJLra/aQg3Fb0M5uFgtzpRMG1c+WhRKZeNq7
9N/kroFvTkjjn6IXPLPcSv8EBmTYRA6unnw3s4H2DNCUtekw6/JGd2KgJ4orf8MA9mXVzArnG8b6
Ug9oVq3YUpGZxQYAXTqX7WsmzHZgMYXYeBX56QvEORTxgZK0jIJEuGOSZiyZuGIuMAH3zcJvDcev
iKl5LzSfE7sGovsCjX1Zvxqbc2SdEad19evv8GjVV4BXHuMppDj6B4EJw2X/5n2vHxBeahmiRB3P
AVYOtspbI7EB0GVyO8JuJJAVw5KopT1A6GtXoJuhgyq+T4vEZG7gjF8oOiITFz1783EokeyFeNGP
wFzb7MLyxxFsiUYFA4gxQdBFeDfy07Se2mGAXHo4Ee7HEiDi+pj0IUfviAOAoyg5UX9Q0X6N2GpR
E8Qo1LdNf8Ln2BqRhz16uBvoiDtDUEfGyCKqeUHjEIUb/jIETL44HfAVlo6WBZPteolmn+XO8Ymr
7WdnDB/LU8nBBZ2Wvz1i60HdsT1pwe47P1tl50t08ySGs3pq5aY02MELzUUO85Tx91pOLI+rVQd8
ocN6RvBhIQVINzTQbNJeS0T54vwGf9lOcXFnBC30O9TC4YyRqrb0KJr4CVCcSourhebiecTSrHOq
WK+mU4DCVw6uBXxBtPoMP03wiuRJHCIk4neQ1NoPYdNc9VhtnUpXrPPeN9eFv5kOo/TnVJZBn+os
Jd3uoxCXnzE3/AdUV5DF0hI5WlJl43zaMU7F+p+v9K+WBXz36F15TuMfbtCOPzC7dxg/4QKXATeF
DAeNVec2KQzUJSf2ieeDQNdPPJ1E/RlCJSoMnIQj5dEb85EjNPqB1AzYRJ5D2mtsBSH8RwRMRgSF
UrANUT0Rbf4v48RhFQ/KvW6y155BbyX8U2QWlpPLtAhOW5br6anh8aUrZleN04Dgod9GbIweRK5f
y1lnRPs14hbg0ySd5WUSdBQvzoGa7ddbf+7NB+ngzGpREsb277yqb4Be5HeofHUpnCevZwZL1MIz
+UAGXwKgd9FWVoIQGC4q3mnFx5Riu1Kd7QYIKBJuXGKRaRw+krBt2oNUch485QNFepVbZW5LkeJD
1pUiF8ntjUfMZEBi5CuBUDDHSLPF/ozKGA9izx70D1Uxzic66XHHuwomn3PuSpPFo7+q7SPVdnlV
3tk9bX94qu0tEu/JQBcVq6YIB29D6eIYl1DRs0a1gfEOQqulnzA22M54usQZs6D7mSTp+WbwdiHs
r6gTfiB5iu18O6BpubZeZJBMZzs/UuxMthVYiGvMWOUcjHMUI+cyvfikMH9LR37ERT3JU6FtgFmq
ioXZp9w7xV7k80pYYUCPbwHDnTa1WcdeRPnDFWg6Y3FlcnUlD8a/yG3t7bNz/cJ65EZSAIltLzT7
JBw2lppI94dCjsmSJxp4+L6QsHKrY7uxPdPTZf+AADTRmgx9kC9DRy4oNpZ8oN2IM8YBE0COK3Cm
fOlJHaQHXHcDTxiFjkDN5iG8ZlNUgn8uh50MIEG3FTUKsHuepG6r3x6JPCD7w8wk5UR2dPmev69t
OdH+uYhKJqjZnMOLEyR7m6FOCUyPxOPXJbqglqyCXqowxs5bKrIZANxnqsSwmXzs8inhQYG9ieSR
Sb6C9VnOQSCdm3y1w++4IauMvxyzqs920Izof0Y39LABrWDgtOgXWjhujz5/ER68EMoB7OYfLrQP
w92po/3Mqmove7M48OLEpFZXjdOt1kNGw8/BPScwYJpXt8WxPiSeDjU7LldHJCEpGGcRfFxgzYrV
aDE2myRCTTJ+hdOp5lBHsYUyBv9jmGkE7ccTltT0nfJT+rHt9sByhgYmaOsYTqLUByrPP45YTZoC
HKvdNnTsPE4wJo7PfHbRBcmt0iGz6JVXU1Wt2d3zvFO8MHHMLaVvI2YlM4+E7PfqUGPC1WIx5AYf
YqjQOCc3fP2YRarTK6hksgH5gEdAAygvT/ZXPFBJDZti07IToTe7dzCqpYm9wzF7yOLMHByXcgak
oXa9VmyNjKaROlo6r6zu1UHTvUGo8oTD15tdv3ruFbRvZS09Gz6OoJmvt2rJGJUgg7m6mQY2FE8s
7KMk5Nw+bl/hlrCK09eKNo7JzKQTPFBtlup4EmP7TKZQio6RVoFuBhJa4VzBnJ920OFj1RvfGteC
akZfZ2/imbpx+X4me3Nv/t1E+R52at6JEczmVyc8Q8i/iXbpYhX1pzLdk9voS/8Ky4RtYeweouWP
WVkTtlWxeu3LrZqKbQMUVZKzT6rLQBJq7ONoTtb5c7W2qgE1550cpsI4mbckLNq+WgKfmKBACwYW
rAmFt5nNxnf8qrHQ2jWOrvyL9JSjQiDsE3KM3V8cH89cMjACViuqn2l5w7zORefDmUb0WE+BFwAJ
p33IvBZZ3v+VIbIxLJliMlXbvteYGwazPEt0qtV09Ii9Q6QeBhHzr5Hk0bj4Jv6PEBbGMzLQcTek
Ay0qv0ovIjD1U2zBuBYG/fjyPYn91fRQkw0a7aOcpzFri0/UVs1iESpe1+ZdsYQ3AwbqeAc7u+Fb
9gm5UNBWXBmXhwUPxogDxaQYX6dh5IVSGS5jhlWrpRNXC/6iqb5YPmnVfEVQlkxyn9YR6aQrRsQp
aaxpf2zKon1RJQbvAR9kX9jaEIaN91RSeyRr5CwqCmfEIs+zX3+VhJVQOq/2IC2vWENVWuHytNrU
gmq2tKJ7+czvAyys/8D7pDv0HjnBkYXHwr1mtRTthr1urJ5pc+Gim9xq2ELexHH8r4Wg1YPKqx4o
6txgGI78NLsExak0AYq+6F/YqK4MPEU+uSNkpWXFFCSevis1QmSp5PFsMtJpBR1Cfd6DE5Ynk/p4
6P9lBgeUmTRp29u/1R04WE0tIPftz/nlE8yKGgmkhLnXD1bTL7MlJm0iIkbvgnrcEfVaDfDxtrMy
flzcPTc65t9Z8GJjVmlf0NQfguZqpLC0Uf7UUb/v06kpxRmM3Wef19lVdgTbFuj7WZKnnhONZMv2
ljlrjJK/JrfIt0IRdINoCn7PmGD3cbcFHATv+ll4B83DZz/+mFeF4XVMbS4aEGPHSbZA54nTr+z6
cYXrTBodysK5WBG6JyNs6ffUKzNt4KAGCpzOcdJ5b3ylrm6qVQNjesq1gnruWVi9uRy0fh1p7TH7
ZTIFLkAXQBSsaUYo/5GgCLDL3xb7k2JS8ui7DLzr6llVIb1JLeB0jiIQB8ufdP8z7rvKizgy6vuV
58O+ByWsAK+zmuQhu13AnyzCtNCsSRyemHl9vudJ/3snDv5XjFNbY0deFb6lnLZ9soh3a5qYkwlo
x/xPhfvlmRKD7Y4R+CKxwlKT5qN0iyByCbTIohjHXUn8c21HfTDWQYz/90yRN84GfB2XSs4j6kdg
8GWWJUZgR/05+mhf1HFLt7HvUrJKSCNSeHQX4J43J6gIttkjCIUPt9CV4xtYzdGVj38+8EiB/3Nb
OPfh68RP1CTjDxzGT79kwQMMQwZgv1FfM5y6vlYIyDO1PPfrRyV9vTNfK9k0ehh6N7OwfroHvD01
iD5g/eA4E76TT6RnrRKbVvneS+ZRB3bqzzqyDwj8IeL0pd+bGbsFcoW6BGxxI51TFAEcHsueyMZx
OgvOE5u0+0H6hKy+/a8SDC00n5CJgpcN3dNalYk15je2KkmKM2oTSthXDr/DW14ocUbijttL2cKU
ZeyvIJoVSX3HBB1QHy8+HO9QXr5a4l8SBul+Ub2rEx6XfP0KG9O2gQN8p1jifRoZdnDkzLqASwml
reMS6ySE3x126yMUk+BxpRPRbHCaSm+OTO/MeShiPzMnqMONS5XQB5XRt4mU3Mmy3Qi2hXE+OZmW
rPA6JgfPfveMyiCy6u3QhnIhO7G+i2lAvH2WuGa+5/D1a9/IlW8EaS0cP6CV/H+gUgCMrLRHcV1w
JPuKnbicsxoPHsJGnvrCh1ihStSyos4LIGOb3ZnWfd1mbtdfRlOaNuU2n6+EyuA1F2Zj0/dxcpiI
kYrbHgzZPM1GA8yzE8/0/HvGURIjzALyhcDphC5hQO+YVHDZl1uZhZDwSLgIIRHzBQQcN6bTytY3
H5N/YTe6X8qwroJu2Nccm4MsZI8KfgRxeGroRijKCrPxl6N9WnWmtPCAJFkhhUtZeQYaAt9OtXdp
wsBVidMxtRqQgI2cpnVDsEvZe7odE5sID0zv/mxP3vQubI058fatCbNn0kh62qRsze4zAuORM5AR
vp5bjkM42uq+iyEgiu0sLv/PxpE99899tqm77Jq0JzSdK3GFhU00c1HW1ED7dsc5yo868OGZg1YT
tf2+b7eZIZtCPaIetomimywp+1dvI/o0tADda0eAHjtP1wytOd49enBZ2QxT5jk1Urxrn6OCcjgV
+ti3a+ELAcIyqlUAHmrLa0WsKgpQgG5h1+hjbn/lOyhCP3epIjGXcN9nYPoiV5PXkIGS/xKFIl5u
IXk2iS1qqgiR/WmHmJDJAD7XvSfJ9xXNBEygjSEDr7C/kOTgCQNVqc9Z9Y5azVssKcb6TL2Gmhfk
C75DaFMlm980wpdhO80togCvnezj8d1EAZt1Ff3QYa6rlm1Jyo5P3Qt+1VY1UDp7zR8lnko0ZBrZ
QNQBp95BXokEmU8Xb8V0gCpSUrGJBVw5pjgjdgTbrxkOiiQBGOL5Rk1g8xpw+Z9BJDFGSs+qq0f0
AAPb+Famv9BCid77xZNPzr3Uy6m4zjn/Q3Fyfdiv4EHZDtnYp/v67pdH4VUni/wGPcO88CVEoYGl
1vEBtPqT2gx7teh3qkRtm46EfTBHWcjT2GVm5k3L6x5g7qiP0o0uO68kb51GGenUk5hfMySAttV/
30pWhG056CrcPmJUmpK+mzO+bLerOLmFsmctw5GE5kU5jR5ht9Z4Qk1WyEVGuRm0/aH8n6COGDtm
TcZGGfz/wCp1q0AmGFcQbatQgiVp43r0uUkDTqjILlDeLCFu8qAOMJMUHOyfBCUmU5OKbs6zWVWc
Jil0J3DgYT+aPK61OP4kKZZSAz1XwXRwcANs+ZFfmuLqAK0umQID+s5JiZOPIFDmRD8lcfZeHPk5
uAWiN9gwDAmLVr9KuGm3CZzwLHyf1NsPyRtG0Tux6M7MhqaxvH3F+pC6C2yqzYKs7gfOqlOyuc+4
GqYI0CDEy7WSNpQu4rOQhlE+Rm+8OvsCpdaNDltbz4i9RMxMCKeMc1tXaUDO5oOQD7XHmaISbhNv
hEb05VF9DiHWbr2uKLmKpVDyeLGcmd0LeP7Qa2TGkxoPkM/4Hn4QudClFzv3tghQ+TQHtEZ/3wPw
tGP0GZwvJpUDb+E8sQHdccp9lqUoVkH1bV5IPt0Mgj6U9pSbz/I/P5OOnJCeFGCOpkhXdEvlhUJV
NssAKdCkmRUc+DeXUWmD2LDwbgWs3LqLd6KOd/hO7o8CyQiu8xt5si5T8V4o4qEd8QYj2e7JiXxj
grEY5nVwEGZgYkzFINWPB/xBjkAlWH7JOar4sZLm97OdpWSXhH5n45ATaKzdf6CWxiajdCE8EeQy
s81c9RERVS2JtKQx8+lxOCQx7afOdY2u09VbkyHBecZQd7TJ0+s5XfkdM0egaOkm4wEPIcilxZTk
OxYpuooxdcRW8kP7kI75rjL+bnSPfaDT/mj/NyOjqc5C+79biJVkZCkO/Rrrp0BWzP1/mOzU3AxU
d4gLgEwyhvIO5PpO1LdF3mrpIGLOpuRdg7kdofRbViarfi0U1szo2CBGNbz/66AElTMcJmbOc9xP
YypTEfUYdfnmUKbZ9E6MJT65D+p0g7FO3VufxohTyExwkF5d/iRGENNZG9Jyn66RgYtGgGb83ZFM
GrI3vB6YNH4h43XlYVYja0vJlrmcxY7EXhWF6WfPpe0/dmVUAMVA0uuw4dEOfS2xFJk6pzUj1JGf
VtzZHAOR7XxXfLehWnbQ7Kg501EE3mfHJqXsr/GDZ0K24L/AjYqqNSMQBPsWvxGjFzgdvHjjb4xq
XmrqKlYwwELeeXRUfAJhrtBIL1SMVJ5H/zfHGnknQvdfB8Uc+liI94WV0YyTOEnPuMoD9Dg5AP6X
OOnfbUaJFnGsW/IaVR+kHgIeUho8kpO2od8FJCpo3u9eSGaBicoTvvL7CcEN7ZiuswtrNQ3RTBZo
9BxutQ9euRQNx9/TVBAsUrNcQXE0zRHWM7BP2i6Xg9X4S2dA3S/Ap7OgLAw7EebLJ3W8uanoAxdo
zJknM4AJhJPseKZuxzgC1yqy05IWRBeiZcSNTg5YOo6YfoAPJE1jx4ldLxYOR2QUKN0ZYJ8rGFfG
QY8w+GUdU4d1xVj97h9iAaZkHX1D0jA3U2OOZh2pZgMUCrjoYW65atzcPb+uYH582QFc14BJusOc
r9CM8GZLcB7RRzb99bggE5SR2IGDu8b5xyoq6/+WScBO9dE49TsJC2AIEut6xfLl5roIwJKGBFmH
iLorLVW/9qn1G49VeiGToo/q4QuR8MD94w7F1TgMBL5A1F+zZXIYu+4tuPEw52C2ZF9MnuKu9sPQ
xebqeY8OvII6GODUxprtzb15vf66Nzcv3FM8BiD5Ssi74W+aEYig5sWm02Fg93/7tjA0hGVzIheC
BA62QRtZJDW5zMtaArL5IsFmcVaG4Av+8OHffdc+i6T3qC9iG2mzEqFlpH3egc2BYRZ9rumcYqgw
mfCx+hWwynbNaVg4IhMQ2Hn3e8Ypsm+wgUamNVFhE8FucAJCWi/a2J3/sUUIhCi+kzJtvxafG4+Z
J7r+8tXec+vghWl3FudtuRyrxSiVf1zYRZARBZXeoMxkyQl4fMYC494UA0JHPW6A6s+0ujKLMr/+
LpnNNqTnOl9prGwVAZTbTYxW5gc6YY8Fxn2kiQax+yr67O/GAeKLZFptGDhekCqAsT/BHn6rX8yZ
ib9UEC6T9ctcmxKUonV6cje4mMNwDhjJ9XEKSt98CmkPyy216BvyC2ShpurFdN4z0+Yd2xodRF0K
V1j7I+3MGSuL/1c338bgIAPWFXehXylEf9WGBJmyQIcKq+l1fWwHm4Go4nRxT/YCJ9W4QspVqRb9
eNXZ3+yKfB76rqayj/RlBiMag5/gWJgDdcdLYjQfwgIsyvtW9Y8zgCokfYs9jI3EsMcDCmjb7J4p
8R68aQcqXbXz2RztWTp9grKEGPAiE7fb0d3eiFoY99jDpYo0c1JnCht3drYmIicNTNJ27fK39PNi
JTv5QR7CxHE+gPpdxcXjox7YnYijGK8x0PpSaxCYxF5NAmS+UONto/azoqsj326AQBHToWFMhxhN
lY/Sq+qpNWYYgOJp6B/e6WzHFq1fnb9adKglWcO12Zj1YSmZ9HvkNeFvpTgo7+Ed/f/sbowph3pK
ZGccTEZQ/rVAkEHx7wb2etOT4ScqbCXN10LtQaczojZ/70b0irAlsJbOog56DLDFzP819aRWQBI2
y+7G9W99Z+FUza6+PhfLmX3YDlOmfh9XrysSOP63KfUNHIGbHr3Qh92eIAMnmAOYMaK4BhCIj4ng
4VAF2ROqst196Cy0cFIjbzQJJjX+lNrW5wekbY0nP8cb1DGT0PSNU/wvTjXS89iqoKP3iwKQUdys
NC8wy+xd1jCryvocSHtCdRoS+dH1Pm8TQ8T3LbBxLu1h5tVLU48iuWkH5t11phvJg7XXqjgLHFxL
q3rakYWmJQDFu9EjW2acHqEMF7lWH0MTxxe+cX9haxjkKPnHgWBzAvpndOMlT1xQFeWqP3foWik8
7v1JJMZohk56Mr1YjznDG5wM1R9mSm2RFFXeb/LuMt0p3bCHnNSzlHQ2WyZ5ccsKRBP3z0uhBuJ4
gpyqzAbYuiBovwz/Z8p8AfXQ+CitASwnOVpAUWLo+abyDGK8SLX82RZj/MUnRr22ND3O+56yLftp
qaapiVQtjZVl50TBnM1xr3q13oKvqS0sQo1OsZmjt+Ah3R5n6q3n1pUW3qbUh9ur7SoQb/UxXIgp
iZlCnrti6wlBL2WhFmvmiP7bhukwoiCvyTVrXo7P9LZEyjwsOb39QBAq0bY1qUzpWyVANMfz/Zs2
xRLFjM7cL73IVW+Ip7P1FFu2e9rR2RqSlpHmhQWns4SPByNQU1iu/BV9INo2eptgD4J4PbqF0UZ8
z/a+ZxkVzGFCbaZqMKW2Ruoxq3JFz0efSO0XvPnZAGTpNcVhn4uf+n7whqLWaKajK2cTfeAXHP6d
Pksdb07WbqMafFcl19WUdsFZ3tWJLTTne/DG0p1Mr2tAHDsQQ691l2ePzF4HKK6msRJpJzA8B+sE
X/N9320HsrxiVmLDgR7igtNMinYU/fSLw6vL7Ih/XLfp9NdAm+8ALGiaNQ+p0XyeNVJgIDwsXREB
Ejp+v7MOBOEUz9Q49T6dSUt3pmS68FvVajD4uapQkcfxqMzcSjGKnxJ9kBrBRsDefiAzcRiFELqP
ggbEU5gNct3LLyQuxh3/MvaZRGA4LRllUH75OvaVKxl+ZbuHLkhdYlz1mESt4qYy+XzUXE7xCRAU
KVxiMZrxwChEk5F/fJPqIwNMZ5gGMeV7l9X3UaqvqCY4uZpNuuZbT3Hv4IkbtJoFHo/Hl2peH1Xq
Oc8iFZz/1whTHvWqAz3LiydPCfyt3mvbdIG4GBYlekbrykSfo/ajqwrHZc1yesCLUmk/0TqAzIhc
PaJfzwg3Oc9lJVs5pL5p9P/ZnhIukF9w9jGUjfc+1Zp5GtVYBT0omFayR5escVeWMlAdx1beyquy
rovP2B9eVlndABvWCynUtuxcuYTl7eIWhK8PUyzZuObKKlB9NmhMpjcZTgG/9n9w502u5kSXsTBX
+Q7Edpr4XCVkx2w3o/vp5Y0hpQq68pSM1pij+zTvfpSsZkZKXiAhLMHgVzpCqjZF6tIdA4FPPNQP
if8uxRHGBxB15z8/e5hNPsptgWSvQ8VICuyBsRjJrZ0smSsNIYdtUGfz9ardcOVRrkqZxlqZK9t8
BYYw/qVCXEoVK1UXLB9btYzZxYGj9jknkL6uLWpiK8ruLs7hjH/ugL9ILvlsNoqnyWz9lduzDbcS
1+fOqGbLkN25bDh433ZhlVIgQVDO+g+dQqvktpDMiSuOXfrbp5JR3PatA29XzaHBayHUViRDmIfk
oBdJGyw3coEXlfKyC1PxzKO2CbvQycwvwgx0PBqcf9aQirbyWtYVGHlTNto+WDkr9V+gnGD67oD7
dpsn85hSRt70Xj0fVMCettOmEMKQg/XWXThPysz1D1ZbJX8eeMuiQNydG0Wyj4eerM4vmx9IrfKI
V4CdFGdg3wLi0XDWtkjpeXgxSJj19zf0aW+fso3cheQk/5ipRR8hZn7o1AQFmubq+JBDg82362l8
yZxZOa/JyvEXDJNVHwJEQU9XtzzRjPHrXvWYIaAgkS9FskOuulSOW+4J8tiSGTojlhWk2jnKVogo
bVHVTf2MHF1OWzD96VyTMImce/qODlSVgjtNz5fSlGvlTMEQmJTIfMtNjrrX1GERZKJte1vSRGop
8ARROc9Ye17R04kh7ihPr6FdvIODBvnxtBIsNkTL0eB3whQA1AvmWPCHPapYQnZiZD5Qtwh+Gps4
aBaOThhGgqO82Pj4UI14cRd1jzJQbnAIme35aUa8vGLAdgSX0xVZtAPBzppUYDXDpTpmvf+igCFt
NOmdaw/9bcYux8qpUA2DCBHcVSjPleJVj2EmT6NDAsw0kLojBvbljSkSkU4kgFdQa4eii4/feBi6
2X5969Wxz73aP/LdoTPPjbMxWwGnz+621HgIay3XpoJ7gks3PKTmGe3EnbDA/hep+tMAU03h36J1
+ptoPO5YrG8Gr7epPL06XfsSPXuT4zgNwVEB0T3MIahY5BhzqgPgCYK7gPxSp1IiCxDdquZ2xM/o
hJ3TkKKJHUIhmQrkNx6i1tZm8a2z53n6yHlAswCcBrMd6gBs1+5j2wLBOtTUGpZ0u4RB44VF9it+
DYOxB/MC08Ke94FFNPkk6Geja+sSkESKHoP2f9wAQNuTpHg4kUi5N//XAaT/pWmIprdWTayBp4mi
68F2V/K4Thm0l9lWt2C3RM/yZZhvkuItI8EJ08V+ohHlOfZNV4PswXdLf1zesXps/J+ikL/FY6DE
v7TcXuHSrqBtoJ1I1NcJR1D8Vz8TNq+yABoDU/4w66X7Iki2I/1+L7WluidCkgrFiyei+I4ceHa9
S7ta5bGKkmYeg9GnDEhDm5x0kC9WbUVAGXJB6Y4iICUdDsh6tsjORD3aRRlD4jsGubi24hOUa4/E
pweJ7CfqfMBqaMTk5QbdUE44xX8Tbf3POvuaQQpfXuS2esnGTVvkhAn2SgZDX67+u/vlt46b1E0D
LxN1jWiaWSmynt6PHagBMuZge/ofKLat2UMflXQpV90paxRLlwH5q7koK7gsYjl8eOBJkMbgJW4Z
beY9DvlH4TymAYs7SaRfZh6EIGtqck3PUWO7TwZVq64xNLoaNh4vDhDQ+ccaPtjQnNLwU1vWewbP
I3CK7QhnuLxDcMCwMU4gqhWhyGje0DIKtqfkD8l1KebTZFtZwMnR1T3nzEZpwJGwUavxW7+aQJZc
ZZaeykC2zSnR0jGugBzIjYwfLPYTqcsNanroYRfBLXVUjPKV7ZtIDidanD0wgsiXBP9wZ86DoyUS
6RgHzFaXSrWW/NnZWxoVOGbqDQI6gJY3G5wCH1btWj8cutVKKhzSyj06tvBAYliRpF1R2u+WiLo2
3Ag1oWJq6mfW4wBEir25tvZGw+C+P/uF9+1JrLdpFJPrDy5Q7SLAUH1yRIeIq9dxrE6AYPypecKp
TktT9kjVfSUAr5adKWFepbm7IBY/K2RCIvSULIOJhB2C6Kbv8I3PxFN8S07gYHo9NE/xahCT+YYF
dCAgBFUx9XwQDw/Po/j4rRnAg0LzWEqo/E+6ZIgbiISaczeICtG+WAtHV8dZG7I45wZAp8Pzq1uw
5s8KRNTrsZ5Tyf9eFrAalPUU8S05c4WaxqPm9Al+s+HPGBkh2fTnvFOSgI6z6Ok3JW1ToQmeqf9J
zZw/IPlAx9nT7ktGZVzvqlsTiqKYKqjyJcofBUSkIpGCLQFt9FBQ8mDMSq/cru0JXR7GUvEsCgc9
1kEBrWwucOzOzOtkzLcDR9OMX4bahg6kP7dMdrFp0WBPeuLiBP8fuBmSmV9+PlOp9zN+T6iqWgXG
z2q90MFkhMEx6IANJ5WpPsQsTh3J9TI5uEAQ4AJGTC3ObkN0ZEojFq5TA6jGw5aBHugGS6gWcy7j
cAXZ0yt7cZSS+B5RhE6TN0cizCanDCfzkIxiS1IdZs4lolTOrf6Ng7D/1VnUdxnZIflxYNXxi3K/
3vyAxzm8AI4aivCUyyvUwvcT/IFmHzjI6rQOH2wJhviQlLCwL45zilVV5OovX2+uMKpwdvL21xo/
0QDjbRg0GrzAEborRF0LjLJq/Dfn3OBKQTLGf/M24SYyBw6s+K1xP3ifW6Pqa6z4r1Ct08okzwyY
hrpyJWDWQc/AC/3Gl+hZswKfCLos3fGp+pnIdmO4SYjvZw6HaJ3mpZ0T4TvbSYD6AfD3LXkvxg7o
L3vBsOXUVL6H0AWF2SPshx8cj2JEcPaYtmPCRKkDy+9wpUKqoiRi1K/m7RwrPELHwpOPubyPO7n0
Banc5aVdqe04i8jbZnJBtZH1zz9vxN5eu3KfOLeO+DqI8R/+F+3T1nFjcfYt5kygzVMPJCG7OWOu
Ws7YQKRt5CP9AfTOisuu6SQMUd1f61amAK53VHUoxCAMD1sSJOBT0jZsoezZhR61/bOGBvZuc1Cq
dmrUMe1nQ+jnhPjV7gjmeemaqVPI5VcJ61P1LRV2+OipEF/zEQOm/5nx4D7QMEEJF5faKK6mkxmR
j42ckwUxX8/jG+11LDzaUdFuzW506Q4MgL++01fZkaphmvoSm6djENmGN8xOGOlnncpPRUD2VXN0
cNdIOzvIs8CRjzY7C6V91R8gpUfqXCv/HTYX1cMtyUiExie/ivIhaOij4rsGfuy9hXAkTt/H+yvm
mNmmuyXD2qMANt/cZsT+8V9TgTLaUe78FGW3mxiMHhFNOIc9g0ENAP1khSU9jyg9MerfQEzFUnZd
bFE0JZj19o0NjTPng+3hm2RdDj30hc9SHYKqUc5mZm+KPhYzcbyv6MDd1gfNvdfGNlrxRiWcq1ML
sgPIMGW7mLrqYjuT9bmHhrD4k4JU+O6zFCmcap71ezhyznO7Y/BZtL2I008MO0fhSPWXfxyronF3
okZocwjydX5DaVGeazsRhehNemOKnYjZMgkNXBci+K+sJC14LpebkPmBKnMH+CtU3kAYwM1/KOyT
VHiGROdvrkGnhm/9lvBHNQHjctwuCFsYVK033TT8dBD1icBULc/gr0NfA1+udi0/CNfUF1zvmGy8
aQN1WjrR0il19hEilYAvcYrwdyfti/T8JxDja5S3BogOaXimfTmjoeS7wRmQ5IPmiavwptu65eHt
40ywKfqxuT8NlClQx8McyR+k+nIiZo9mTLCt8kFIZdmdLo+X1C7e0TmiLAZJCDNoxP052I+v4hPt
pvVjgyokxjLkshT52rYo6AjyTzI88njz639ALIriQ/MggAGS3yNJPCK5Xt9YpT1ssg0M9G3YNzFU
lQt8frSMOGbhB9axOwPtlgGHRPscJ6ytMP53hc3cxzpy4IszMpu9CGQjOGtIW2dfE0t2PxN2wxgE
d0U89pNiieS9NbuHaVB5SiD0UZhDEql/LMevP1xq+yDfUfmxdcJYTRYqzGeptfSJ4htyIVn2GT1F
FVfLkhSuh/joiEaWBXgodjtFgSNA14Q3bugEWjLvEic7EaBceJjWXTZnarq9rgxI5HA8eX6h2341
WIL/9aEB45qpk7dENqpLYfmwnQ7uBvrXUDOXxtZoHhBAhP2dDiIZZ4+JqSyKbnvxtLFwt5xLTTFG
/uejzIyS0OzS9/EefACVB8GdisqPYmRr0hPton/wM0m1os6BWO7jfTGIWljFf5KB5VHz2KaGxUvs
eZgiOpmgrjwLjUangBHGznYUI9vgRs6SuGOEVzWzZuxqDwLEeguHwLxqrBNFUJ1wSKBdfteE9MRu
9UbhZL4WwlGKk8+8LSRy9BxcFMkO+rLQ4udHx5sTuu5tJ+yYgxVT5e/1DXFMhb3DtW8JY/CNhPHI
90f1KTFZRUAcLfOPBc5fTw18KwjZc5B4JzUgblT3la7GCU16ReLLx8p4eeXanE6HL4EWjlba9yGD
toW2HlRo34IYkOuvMxIWQ8X9wOselOvC0Ayb9VM1B7aOecs87UwBx1RdRTnFlwSJxF66Y+UJX0+s
z5DUEIYilnA3efCjj/4xcCgppmCzj98PfdZLE9Rh1YkEWnMRg4DYedjkrEFaZRInM/nR0r/JMEnX
lbIiGmVAv+Umoi9YXiiq7ZMO9smoD1E7EIGnVT6aztaiD6zPcUdunSv5aLcXyVkj9ma0J4JVFP96
IwDBdoJWLc1VHGkZqt672137qZLF7Ls9mL+VzpLjXA5c2TxAvt5NNxFedijgEADd++9YAUdzf39C
+POLqXOWdUabjVCFhwYLIDJLj6duZMJIauFaCSrhUydXVE5b9gwINWBQhjCMsT+7H8kuWXbNSnhK
m1e0li8twTHwl3Jcg6lGcPQ9qsvK0BPuhaGwGDde/jBxo8qNS6A2Sof5pAbvfT6vrMfO+uXP+n5a
2J8xo7yYzrWqBr04lYsif+lR6BoFMH2yeFdzUHacMiQGjh3pnzo5pIlceuTmG1QFc8fYAUcbcw9a
8LbhgA96mKHojPzXhDRdqW9AsiWEoRJXl2JHHmi+IfRIzAfcJ0vwU1HCSMzU6hOQ4n9D7DCUKgrt
ORq/R/29EJCxjyCtYgPzuplzuXdooBS3lWRF0XiqFGHOKxAy6+MYqRysffKUh9Nucka1PESw47xt
KLuGjjsvEYuUorM1KWJvFR1t6teruwb7AtSuvGJKpN50076NviSgBrgugavanNIywq2sfcTe5bwl
K9rkDwc1DHxOBLaZ1Bl5h9u7p5lOYDiGaDhkqZSNaqHIkaS1K5YLN7WfmMyPjuUE/OH6KPkwLauK
CKDAcj2JXNgD8dGyEG2aS8DtbAgWlwR3SMemMIxeF6A8o/7UjXtYKUM/rQYByrxjZtjxjYymQkps
SLoOqneZ/rDYez9y9o2hahl52mK7T1yWM3Dzf15XKfiKeZyhvbnXHNrK1wNASYJUKAaK8b9/LhA/
TX/jQsd/ED/FZtErdAVCxnqn3gkFtRpv//IflZAgeqJIJy1EfMtTfOBDkzI7qBi1uB/0taHWrt2U
hxucRYLVIndQlgl5ii0rZbSWuJzSE3pUIBOG5Lu2sb9iCZhzP/PHyWVPvnNc0VFD/QKxeLGavM/p
skqnk+hEKq31ARWEohtJBahvdIVdkdQO9aIOoGEr2Oz41OGD+dXfxcsDMdqbHZtwPEk+OV0lnDLb
PlGUpgySgVVygR1zDfPvx4MeiSV9MHHuSSy0ud1JVlJJrlKsxP83gQQNku+aNW21Ahi3vfIsIv8S
rtNleunPqlF+ruhaled0hNwmOUVRJeFDZgmwrmX9OtvCEeFoDzIehmKElHvFUWDP9SOHDFVdiCAF
7frH9cIpBptLONU83CIgD1Gq0Y/oKEPG6jQT10IWIRxWyaWVJWZttD/cTwaZapnFktj6fGRrxobg
h/NAkE8hBfnitJWspE+b6uivWSWoskdYlcvb4GE0eF9nOzuJ7bcIXXlP5BrV2EpBOc8R5uGxqNZP
8NGTccJttt/pie51xCt3/HUwJmveDr/jHWDAslg59GIA8q4IifrBxpPatrsyqJX0YLxY0lbVl6Rg
bzmz8cOJJyUYfJkrKw9OC0aJSWiFRgeJRPYtdNWwFo/I51L573e7cI06wzDkEVFTqWzVAsqoGVPc
QDjy8OFjy1NIWnhveqkgfA6AR3AOFWEwVJ0v1+nEV5FrUEdk2GdXYUxr3KPkaW+mvp5WfC0zdqgW
GpxqnzMrc8Y9WrYuLMYAXIZBl8r0gEisN1UG4FV5T/XxXH42cj0TDuQWhjXgsJofRjdZ4FrwfrcE
NdBCTDlIlvV5gkOPrWB1surxra85YocvDVXJCyXmwlzUnnM4e4jT9obQqAwZjA8Gpx4Q3Mz+u/ee
oWx1U4FUvY1lGMp8B3ldW4fSXVFvcPejMrKKwgb9yUURSFyDiUTfhi/3k046yM+Ekx8nAC/gD8v/
ksEXlDqajHu5EFuJ6jaCF03qZFzsF13K/2LIymt1oXfx55PUuRVo5gkO3+JIHsiLrRatDyj1D0s2
IybyZv366e2KCGHaeW3PU3/WuvUwiD9VbEoAiO2AxjdgwLk6WYyeW3v87fqbODJcTuwm47J+vEpO
wIF2bK+GU68YHOtUZqWwmrRx74DEByA6FblPwN1oyfgRfwomcyDlSDRSMV6bVz1dzNGwLX9ODnUX
ZTAKY5OI/E/lzw6/PJBGcrXA9fZ/IW62VL9oK+4WSUw5bGD5XNjENzjvYXWDTTDaftUg+ytPRZ7a
vTacGFM2tKfx/hdqRHcwf7yUU2zuaZfAP0oAg3KxgTx9keO6n3evLKPF/fYWKPMld6Id0rVdiV/d
WDzRCFOiSbsaoB8NageuSDo2NMwSRPpFxCBUIHsMOPaAILDvJ6rVy3kaIbq6ehIGjoBvof98xPrH
J6ABmQIFitbNmxUdsf73d9YbrWW1h2Q7NM5Am/FzpQU2KmM5exz7HVEoEwIxW+dyIqGhuysQKQxE
i+DM2gaerUMcSC2IB3GM0HepgOgqEp7aXKpF5X5ngl/RHOuBudiSuaV4VoP7odSj8THCUayAJAps
UK3hIEAFQrUtAQOZqe75MWVZJcyNIvKWy5lWc4GwkWuZoQ/Lu0EKJMEnSu4JsgF58D4MVB50ruQb
0OhzKJlMzGP0Cv8WF5MhDmIkkcQgh+8cqDhWAqq5PHR4dp3ooO9qSifM8k6CASb8fiaZ60y/9CGi
JqRfqFNHJA0i2V2V9dyTUWT+bl0hNX9YBkKIMUVL0LZiQsjZ1htvCSq3fbX7v4Wj1HeBYOg6uB71
O72VSstqdWEh1+BCaQjRoFnDuLcJQV0ZLQ0RhHU5AOvn2bq+7b5U7Aq0CJ7qPUJk4w+NoP5demkw
V9IeGW9OITOZ9S6WOgJ2+cSzYT225wu2ZsQaW58c5sJHf8OjoYQl8UVEdGVMKW8w2a2+ZWfDxBg6
vmRdREIykbRvytIb49zmBOeiMBYMeJlF+gBjWIzsohD/coYsldW7UtCvRhEW4w81drHGn0v1Ww+U
LKrI7ezf1HjP69jT0Jv1BioJ+7Ni3CYaUnlZiPfb2XpumB3p0oN8Y1Kt70P8eHNcEHIgyxfvtPyB
B7c2Wedd1Whbry8lu1zMIffV8WebBq2PHRrGIG5bTzJCEJ7blzN07+U8B6blxSuNNw904zV7TARo
W1E8HrfDcx0FaBNYcpyfCrI7mbCqMuDsI3i6eAQ31ZrXt94Dkxiyvq/SZWhGcLZx9vM+Vzu+y9DX
lfsLlFF6PG7spZ2N8g9paWuExB+zd7bpmNSIAGUlWVjpNBa/FShn1/Ot7mR5dsyq6OGxlsJObfr4
mMSPs6ou4Tw7LFedrf0NbAe8B6dsLgOkg5kLMxp2CQIQTyAytzSoLzWAr7YxToTH1m4f/FbSXI3u
ocjr54MeSHkzLEFtBm6VTDhB/zo+CwmGlp41TlxxEllMRZDNhYyQNyVlTZbEasgKR/jknzXkRt1g
ikoC9jj1IsEXwE/oGNaTpBpmSpEoodwrzL1UDsCJurYqYbGcwwJhuQPCooaJVIaZJAp1nKteDsw+
hZSeaYXZAc5tx9L4fL1GWdwkdNTzCaedysQZy9D5W+JZ13CZSliER2U4zYoSQ0pC2wPoR1yENifh
ttG4aCQwW7xp0QWGxgQy1RghaXkT1YNSLTTPPdlcSFmNmra4KEZUm+TnBrQk8F24Qn3WQMu9pUv2
knarS7WttZICQTRKuDW6/8LoC7XDn8ULxo7DwDB725M2cgKCdUMEFVSLEEPFLJC1mVYGyM52Ek/Z
8Yi3PxHrN0ZZkTKYp1wKM1was8PaflsypWf8gfbMcXUTbwhSajeUyerAW5jnjuruFBuc93h9aQCM
HRJs71DJ/uImKQK4vNZd/DID81XR4qkBAgHAFPIvw353CsGb0++vxtdLmUIln62WKo+uDvBaZcto
T4WXGZ1F6MB+39w0Zc0n17ioUF8RljDhs7EFafm/j02UOnyM0DxkVqauDbMMXF5XQCpbE7KKgniK
7iJ9cbRyreqMcg20rz0ZKvXa7P3cgDJEyikgbNTmj2Pb8AlYnGlSLHM4vQBYkZOKevxED6+MJ7j5
slIvDjBR7yuGxPIRwbiXT/f3upMT8+9D9/fF5KA42VV631JMaXYvyW6XjbvZ5zWZc5YZ7DoLyCxK
rGckBxwd5FymPCAOO25WklUgyZPGcg0d4okLspTbocevhd1fpx1XOrhA3rOX0vfhdse78FQHzqw6
4gYwNbNXZGUw5ZZAZlJhqIviLM2AVBThQ/0casowqnOhDVTbfs30jJKABNLEdp60tYlnNaNnXeXl
2SSwjUlfUSac5obF2sQ4k+Uszj6MhcVzvpRI9AwYTPTFPfNK4Qed7b4LzcvrfWQV8r/Ny/h4ATto
Z0m1LoEjL3MZ1ewKlfFrwp1r0Y2ECP2I8IDRiJOY36lpOWX4+U/5vq/KzsHV/JSlyagEhS9oDlwz
x9wcqJTeA4wot91bkigptE3EcqVqKUkQTXi1KaSHGiieiaGHTAN5/mYzOj2BWPlWNUqUMUPe/mJs
HMo29YHhMxF0nGPSkay/IafxopYoWe1HtCWPQpImjSqox0+jJNFx5esk6xOaJvfQmjNpADzOjcTb
SfX1ubMYFjrkxOdCqbl/t/taLF5nc80uwoIMu45ftcaL1tStcEUoHjpdOI0nQogte2FrWVcKJrZg
P4u8BCk45aJbPrTGP+8SXdzdwxBRwr8o5MhOUMMkKzKpGRXdIaUBkzv3LLadKTLgMZ6FzSFbNGsT
KmnqsYirC3M13BHhjRmbihTgqNuTXLcg7HBxY249mFGkyeepISn5wIPMOa6J6miRCi12VZ8V3b0c
5LWZAeoCkrg44n+8GZ6TxtewWRehNZFTy/hXiy696jQTJZukHIcANG8/zxCtY0B9OX6vPvzcc6DT
94ktVktw/MhPohTelKmze1AB7A75AzyDGpzUkOadEgMkuKEWTBM1jtsvm1pgHpRdiDsqdtUUjc1E
ql/zgDoRbnEMME24usFjcAdrANgFD65OtpQRy+WXE4bPODhFHRkrJjtT/PrHYTdfX9uKUmSw1W5V
i3aEiy79wWOhVS8v3CDcW9i/r+lZMdE2ezDQd1vubbooHpPmN9PKq3b2Ue1bv2j0M5ZH7E2OfdLe
1GPCBnGd24glB3WvALCRGV1lm3rkmIF8/u/TypKGMJBKeiu7dOicRY1I11/n9XCWeW0SCpUoQZEu
Mq9FfwwlBFqdtZwpSTBQRY1d2Oi2BiVZV5MspT35gf5jtcW7fbsGNYoN7lCqRM8GR+YGXMSpRSwY
G4Ue4NsB6GD9ZBbqLHkaz4KIjgup+1BjzMA6cCu74plh0oBshLtcZHq0T0S5n0voDG1GeKFmCQu8
A7rt3oT6si33n8cbARJTdM+rNSOmq91+/XKfhSFXw5XeUQA/6JcbX0Ylr7VlK4sPo6LCHOpcQSoj
5zqi8apnbVLxhcPrngbDomXtZtqqwqNn3BBye8P1BL+qJo7u3n9jMA3qoWNb8v9QwLPa9M+RytTQ
8M8Z6QBWzO8q9qDx6P1c0cFgFkhYsbbDWobts4KVptf/GoziscC3OgtWMnKobPczXLQcy1avU6sb
Kzjo4bX+1+XrzP8paCvIT20o5J1i7Od1cYBNMRp3akrI+f4FminmJMhVBlrsiR/neXOkYgPLYk4H
p84URW7C6u4PXrau/8HNKjxtwxCNGGC3MHGT7muoGnte7WjsPnOLFJ01IrvrTax2nYqVMPVfP70t
3kBjc8v9uw78BsmzfQwGP//cMMdV8EDsqzTnLL8jPJ6mmAJua6Hxx3QAgMm3vjbzRGGKsGMqtaSP
pmRLYvI6ADKXPoBpEvEBWdM/Eg6RhMxeiNvx1A9TCLK9Ob+jLp7vChmwG4uIRZKeKgHGE06z9Rkl
FF2bqYGFKsqFOmaTi4EoRvWtMpInt2coYvks2CC82X4wrJd4jN7gYj2R+mzWGAsbNFInqQytOLFf
H7lHdaxCeDDIQ+imSl1K1DndeatfcnptZtFTtgAWp1Egps6rJjwR5BvCUqvapDM10lQfJM6pOL6S
K8BCcd83q3pLnP97GCqErDSXYTR6zw9Exjof7GWWxScUUIeH/0bK0sNszYbqOTf2+XrVhKlby+/h
bhn6ZwvEWZw25IYqKgAx0CaECKF+FHqabTE8LxkbRjPrMb1Wt3ghl87B9UL9509DVnm4nYMTD9d8
ICcnFlHVbSSDzwUiFpyBx/tl2d0OdVs2rWp4D1kBUsMTFbXKcFUf3lTiUdAW4vEVRQLs7l7gje3F
/kXvelZ514lFZefXClFQBxPRRlUGoBcTMPAVkVH2rCh5N9VcNTIw++1EMibb0s9ZDumb9f4KOEaC
n/OWkdrFVEF+mTZBa5U+cPZG56Frw1ebE72AEnBTBzVE9deDho2+dfHyoLBsqb/8ZHVHsX6cLYQn
ysjjKxMDffzzHH9V9Rby0KL053ESqrR3DCKrmY7PRF7UGRd7zqm2W/wkJc6iGX8HWOmW5fbDWT0x
F5xkoWiRLDpZdpf1FkuXgI/8jRft+kIHRPzq3ah3LPn2y2xlSMUXssgOilw6NtJWHMBFJcdWsbHG
poxLz76vNlvhm3ZSFKH0aqhaIRxo+qTcsY2xP/iSGxCG94k76kYPShp+zbI3KDFh5AHB1reUpOv5
n8a3P1Z35xt5wVStSBNgoshRW7i+vXJRQqQ4ebV24hLjxTrkHyFY7CyDGtKNM0/9lTZBvDqha+zv
60jhgEqeLJa9R8lLzTjcmLlY4Z0atkuwkxcrTrzfMwxukXf+u0fSzBucIL25CimYPQSLXvEyru0S
UoWTs8tt5rjFRyg9DWgGPqiM9/hUCl9MGOgzWhMSDy0crYrGrLawFbAvckZ79PKXyJJABd/sr/e7
qFad/Z/96ZU9h/NzjTYPHPH0+KT3avTJXN5jbj+Yeuq9ElSmz9lFMLxUDlRyRFLyBmbsfjtpWz1L
Cin95yYs7VXrYzXIn9aSzxy5Afs0QlrGDTO0WQ1TYhp3E0UhxT3nRIQibbu++dDJXluRG1LoAUG4
COTFzTvVXTjeNX/C8XS3I7RRdMJWVX1BenbxWqH6m0LVcPgco9GZRXZEUMBaoBDgOKkJThuyu1Kq
w17u2K3c/Eg91isd7QzjnH2aqiFhXOXrnNy0kdRuXc0CWlIcJVNXwRchea9XvhwGzsO6pIh036dt
cisKq79Hr25Ok06eIA0d23BzW/n9QoGv2hHyUNm22+Bc6BCgtE/u/CO3COURoNvrb0EoRdujSq1h
B+ipPIHCfGqcJLyEUFljWXCdISM7wBEVY719EAy2yZ2aYDbrMdoSXsVdVOCnu0mFXESZxE6c8Pzg
MOJmS7QaCqQWjqyYMVpM4CJOfuvG930ImfM1j9uT6hoZV4EPJtAzjK3o118vnPDvO0m5mi8EcxGd
a+Q/Wwb6cshm49u6IiS/LizR4JKfx8SCgrnhjopy/PfAZdxgc7qc/Efix4IsxhB6aQJzJ59PopQj
fZ4t6MsBvosfTLGIL4sBNn2P+2NPceCfG1GD3nXrbSz2T3c8+SkUTN7Me7St2I6HYWWXwx5Nk0xv
aeZG7UcDCm0nYE4WZJQr1U0hEsSTlWRGp/ov5Wgm5vnNh0+DniqDazhWMvP9Gv6GV6JBLm5TvEMW
IrfUVPgfN+AXxOiz7dXRytTGs5zTuvvCMCWKlN9irecBsJr2ABpTtY2QEJOEVL39tD1ZLgirc1V0
942r5hCgSWbDY/V7MMOXUh+NXIdqbCF2glLzZDQP62IVfXkLcnPBgXprvQsAGVWjNOJ0AuMiZXyn
Z4vyztAkUrGnBS0N69+kYfE8RC3qeXb+0fJZHFFqGz6ZalUXdrZHaAzm/XCl+yJvuO9/JXtRllFH
CglhRwWdBairaov0GCylH/bAKJ9qF7KCKhnjDaOUO8CUNPiC+9fLXkY4nIBDrV9gRs8eRrLuK8Yj
mBEQApxXyAtSEpBu3AydJe0T36N4dD82vZKLr23YnPz/0r8TgyZkU8t7gK5bbc/X7icQKvN+DzFV
M1T1qJ8Tqiqa39uapAidHVLEzjM3grdB+sSnisjevOZMp8nk8uKKC3ALEWIEvvPCJenk51v1xYlz
fC7hytJvqcUJwyOuCXQeZIC4XL2md0Pv4a3kYRjB2qawEyXYNXAviiCRNe9oiy38Q7lIvAs0ILTS
wSMuWY7mI52U1BEhb/XgwQnBEr/MBc4LVcmmDUCKDWFXZMZOsnyrhfZOdZFrKgRA3FBIVO1P13gQ
EyvfwAM2T1ah+/C0iQkBn+Ag63Fk7LC/gkbIzHrqTmVu0AETEsr994U7cs4ct1FdkVqlAIyE0ZbH
9O0ofFyJfeLM2VHf6RR+X4gIR81cObr11LFxEtDxaDH+t7dgPIn8qqJut5fIltvIQ6UHcgbWR6zT
DZJZT0+j73V4V0k6YgI0mM4aeFqNLffcBF5wl0s5M3/ZIh6RJbxXOa+qvjtnPNJXqzK420u75gpm
a2qNqzyRyuiJ0F2Ep/CKCNTH87S+8TL5QTK3KDvPGfIVTWNeYR0ZB+FdhFLjspYiBU47QgCRR2Mn
QDGKt9RzAIQ2HA/gVLkxVi5wksUO85ggdoiZ2/tSifrO69/ClEmfxDO+AUnYQ9yuwS0pxHHBJxj6
zQlSdwCaBAk60aRZTHWJCf9HT74Xw0o+pYRvxgr3J5g4BdyfCIFyTIPv4e02o0AxBvLkRUQGAkWm
Q1cpylvfYp0DJ1El8pDYZomwbuyJyBN1ee18cQZIlTzJnlVQo4p9sUMFl9rdhXmgs3dTlFTinLB4
8qoRXPwmIYtueEP2mdTZbPRY0xyLpZGgrJFecCOtF3aMhvSOan01DZ07Jxn9iU4+gzSyraPKN/4a
DK9jEdck+Lu02+vpUmwBDgQj6DtshDfgSA75vBAp0fUjiDTDmbAUtw1Tfkg3I1+wAV0Kd0YJgqME
hevXQlo5zP3Ed9ZwH4+Qk6ku69xJQi4nym6l7nMgukZUgh3yr0JcODOYXOoMg0mh2rdfZAZPoN4j
62HNmYAhFfkuLLuWWmuOvaLrlZ3frrXWHeGwAX+8tqX/4zzZJad+6jQJpayIUPQ/t+fmKgc1/yMB
GIDcYElfOH9+2nksq/JKBIno1SZT1YWRXKQeNbol9cCTgKgx6Kz6ZkGVpF9pzSujW0jF6EmyuHFE
0HYjyMV8xPiCCL95qxLqWdA3N0xongOAHuNq03pBnkHuJl6C3Y9ic94+bM0VruU5cTnewar3VMid
mN7COnAwuZKYsk3xHbBgXtOy8UFZa8MUMqFkLKYK0OQNc/CmXCpYCQndQiCmkCFnBsMt5LcNXBS8
1TWe37EQxsKrIwVsuKeUNQh3FtHdCmEpXkFd9RJ+cEy2MAzmwLzBKRvXw0WgBjUaQh44keOpUsB+
FxU3j1b93pQ53h93HrcFshIxz7AZG5S3g9MI87a+oFMnGkkPbDaNUo6+W5sKhaesTWRVho2/49xp
yfwALi4FNBavimudIl7mNw/4FFPx6ybTyxD10rWtVczsxMjj1m+NpyZixj4xQG0G5aw2OLGP3899
RlNTFOeRBaimWua+Y9TbYAUuYJ8/2xoTII5MDMM3dEZx49s3ZHsTVj6iZgctQ6G74GJorZTaNzYa
X8Jm4WV2Y8qsKZu09s+JZrL0Zn4h2riMbAVg+XfY2ggIV0YrsCSNbSXynrFvVmLCoc+3uQ5L1QsO
k+ZKCluvQ9ekLKOi+SbIxc4GwO+1dLfeDDlHmjEG0qQ/BHH0cON5n/4rZ6tKIRz876gUkekfETyk
Zw/q6Z8I3rY34+xBnIC/WjFRKO+DhGpMLgTGerOl2jNBEQz5nANc2oH1YlnxZv6uqU9F0VERfXgX
pUdNiWdwkSXgDXfVg2P60KJET4O4CGQ8XderHCHA6Zon6/mvBEE1E0dOSPAJfo1WhDxY02slR6m2
HbqHsvEe8m4mTk9knTUNUkzwey82E/KnjxrGo+QO0YNEdMwrftATS6pbzVK3llGEBwVimyvkwk/x
SYlEz74Ac+9GqdRgDuzScXwWBBQOZkUq8d7aszvs4lc8t8heDLyfhis5thXLk5KlYGjrkLyEFYJm
cezCs+6fh9Qo+7rWwgz34iTNgAmpkDOfFATRYGKyLL7SyJNVrdfDzR3QWPQsSixXx4/w86J5YAc3
MWpCCYCPV8U9AoVMNsK3A8/KzoKiu+ILhUgeFvJOWl12lnuRZ3VgLotilCmEJXT+0sCMk7wiV9Md
GqrIYGK1e8/YMq7Rg/2ozKF7GJVCps/n7zGKKTqvzj4uPJSoqm9HY23bjVNbs3UH4fxa8NLFxasg
INfc/jTSVZXtqrfxtYMIO1W5iQGWyvmbENaTHfxy80U03QBrHZ8Rtf4/+MYXUl9ZqGGmlAys/54X
Ic3k4EbXTpQRDFP+uM5nWgfktZlmHsQcIyFX4x7ASeJVlaI6uIhdQOKEVuZL4JbgwBPQ1JcQTm1c
9+4eubKbXRDktW/h/noPp1f1tkm/EWoHHfaTgv47ScbSKwr8jV2lgg5+aqHtefO8LgIYXaZmEwpF
c8WGeSWr0OzcvnVlk84s9DVjWzieg4nCel8LkA0Zag8xymxWZN7YYTo+Pvn75BKuXvMNjYiG9TGK
KozdJkukbWvvv/aqTMn/ivjBDFbXr3U//0TB5WcS98qLexrP6PhRJd3fqJu97yXve3Y4KtgOWJ/8
jJhgXfCQA1pr/tcxRyum5GPzvYCr57osasjpspmbv5tMevVonZySV4gSw11GQv/R+WTQXd0xW3gY
NwbAFiCO0q1GI22667AtQT8K8l76uRD5CDUnmtVV+zn4AfQOdh1KVFi2s3Ef878/kP/jtYrePI6I
GOsq2R/vQ/hI2hhACxWvj7a9xpAZ0wd7htw1laBsR/mXGaRO4MwcmXAg4ku8+K1SNDcQel0mnzmU
CsznrsUyOFlT92OFK3Ooy33lXuTQZA3yh371zbfFzCp1BYYGwJDuqzOQD3UnV187KAb/OcP2XwkI
3jqyg9XY9mce6iYWwzTm2/vyI4+aLUwoW/gu/LrKOyrZr0WGT2OR+2wboK5QqxGx2p2NihATU28j
f8Z0rUl5axKMfqSC1q2Q7G1jsi8xQWVIbwYkFitvbQUkxLrqjhPpTkQLL0F3vVN73X+4LJIa9jej
CtYvkwMS12/8ee9mEBnWv5I3wfE8j9PYFHws9Bde+uJkkPOfVsxzu8uOERbC/LNAKw/4R2YX1+wJ
Uqfm4nZ9+g7FcUbtCoXCH+cGaHDcAupJZ9sFywMD6WqxhuV+bUt4kEsqYQbzcOIEm50ByQME5cpc
6myki7XG9UFopME4vDGmgFZpD+hPwXtVq4Xu4KXnYoKuKWJYFRtxJP0h1R2I8g936oOMal9OX4mW
oV9B5KLD1OmrNSUVpFHTquAyQR2Sw6tqQxFq7sm0Fn5UWHu2ywv0UT96A9vH6Qcix8X/B7JRbqtb
NHYQ9Vnzcg83l/5urBX7JiZoAEOLV57jdQKmht6sSxWCGuPTQ4viBiea4mYr0tj3i0CGjuNi+K66
ApafoP5lb54kNQF8DVLLmcAG7JhGHxbmF8X52/q9v98ExoNIeWyOof+H507KMViazX6SKuiqTAT3
Y64XaO/c9SGtZDT3yL8ycaDEYc5wridfUBbJf3adDfp1cugHnMmGZrwxjrBEKUywoMT7BaJkIVTB
+QNWEppV+EosWpOnkaovvkRjUvdb0luED3yC7BTiDjBfuc++CHmWxi2K82xXciyYS6AVvVYH5opX
HXcF9q4Pb3MTKdNt8+Cp0sCTm8jtfln1GBYHr8q/Uh0ldJRu3tbz6WxrB3kodIskzGIYmmeJW7nn
4K4fMR3+DigI8eZ8ShkDGu9oz2K5CenFNPFoL6WXnvnE9pn9cZPlv1bzFEhV6UnUyWeQt5LKTsaS
f+VwhY4c44RdAjGOe/oBxDLYRtdHj0DBW0xn8PjjiGNml2cDvGnVOZ+DyMwAAH8IiVLUaBDaksi3
AzH1Qed4ZPzUlP+S9pn+xLiaH+pveRLo/Q2CgFeSU+r4WlMaEQzOkhQhz2IQSl/98XfYfmZicGTJ
o3Umjcjw09sAa9Ob9RKpSMRRu9W2IyuhegwvJU+D2tRxQTr/Q9oSav5qjwFJKKjZfw0SUZgrjp+d
j+qgVRCNcwPsVFArGFPgYBRIqXlCfxB0emZyg+SL9j4iXx7WtvK+Dw5Y/1zjgRkc+xib7wE0fS9N
tBx9q6As2LpkV8jFxS775K6oPxARg6Cg0R2ukk8uYpSACzrxPvQWRZj+NfCOXAPxR9OoLj23i0Id
xNM6c+YBTE5ZBn/tU5YmfM6RnEEDn3fgMJ3sux/pYZNPycvYrVjuKnEnIy5ltdOZdSx8VtPGxLpI
YjFAi3nupVn5Z2kWeFk2FC459ndS9er0m9s3bqPUa5hR4J0/X7fYL24Jtp/Aq969xiknEGvZUOO7
V3+QIYgM6uMTCmH+lwHDPrX4oJLxZJl0rA+TBiDAespZGO35E6CbM2NTmTlzmyPyicMAWQB5R2Z3
Lg1i8fXr6nzHF6C5R1c7PDDo6i4qv3qq378RLllPxYhlfzugsLgm1ltX/Fey+uh3LmiYPj5/cZTb
oCvYqej/Jr5XZUGD3sAiORZTzBZn7E4DJ2BH0hohJUt4d+vENNnRS/CdWhqJ0psWAE4tyz9vSqQs
zTI5Y1CQRD4wcx+LigMx1lOfRCoV/ZUFWUQsGr0UhjDMFrnnxB3ICjntPL16tuUeZKpu0F5i7lcC
7owGmUHtMxxFXsqT1roBcS6pf4w80p5rWdDwPEnwPnBippKbCFBeN0Em3qC1Hiy20tmaww9jSGNb
Hq1K6ZXcNTzg33NWHBqHQyJ+8G0Nsf/UWcUhKFU3m1YO1qFXe5pxP+loPkh/qk4i2pA5c99q7zos
tFpX0q0h4yukYSNnLCuUv0pDx1sXT1wPvdNW8CpDfFLSQTVi1qhj4WobLBtpDvTjV7+XVmUXnNcP
co4H8HyeNg/QCJATwAgQOLAeYd894zyRuS3pE2tjGYmhCDiGkQeYdmOfPsgWEOCBdrBT1KQ0TPxp
093Xj920ZTmjYOZ/5aA0aDeFokIJYoXZmxKKgh9AhifMlCasg9H4XcNM/sEvDSLMSwu/lMeE1sqh
NXir4L2QzKczCSWoVUGK0oy7HcqASFBj/8zxiYQNR32VKN3DNabyHb47xyDDGc+lMm8OzH/ppale
GHj5JanAVETiLuE0OEFw2Zfwpq/bgrN9ne5P8yUjTyvXSgPLqy51juSixnPMzwt77e4OyoQ0XfGP
qhCxXe/NgepUzehdwqGjAxCM68IjpY50tPdH9HFAUzSEmx/y3Mld1D04gHvETjdBkOzC0c9u/px5
kBIZFUzoNHYSgWrRHQ5KZYF050xHiWFt4NjltzgOacpsoi3MVO4EKVIomWw7gfV7xCKrMdUa/Seq
rzuI+8OhlZOpIXl9BbVSlIPZZ/a0brCo8UmIFDpmw9g7/sF5EIcISnXyqDoeGG/hL0v4PY1M4X6P
YTFZC/sr5nWj+VGqkW5aHEyB7NSGpVZC0lCn8TelhI2rcU+cqWNYA7Fnm7Jttw8et2wfoQKr/Ke/
/rpOmcjEfnBXK86vwYQDY4fXte8aeYLRuIHa2wJvUfrhRa33gySlZy3kq17+37YGER5HRwYThz+6
czendg5ev5lJmeXPRz5UFWCwKEf2oSNV67rTgZUqG8qShontB5oru4C2JxozQ1ZmdxwXl+lHy0VS
5BJA276iz/Ho9rz8mHVXllYXfNiARg7IwgbvwMR2Jp9BYi86LzSBXSx6flQUVBV4K+6yVK5T5/0G
JeJEh5xFeidiEF6WaVO0joEz1Bm1TbXabIYRR2gXGqOwtPMTmrd3OZh9Gs+m/B5l0Qtg/vbnFAjs
DWRnf7cm4q26hjVi22/tFdcbbPYKZ9fMfw+La9TiA28Pqqt5YUZzRe/lRN0a8A86ZuC3uu2Yq62X
mDGkTaH9mPgF5mc8gvFdGsOXuxoFr846MtWaiDG3ZE79dC/ofj+XbobuWnZhd41J2/DhkAekMYUe
y/NCR841KMPxT8uDjtaAvbZv5RKQIcDyT3MB+iQAVtV8nzxERqd+VfuKEks4pW2aPr68CfmigEKy
XC6iPOec20FyEvgAKCU1T6r9J7ESnCrRM4gQxvftw6AYRiMvl4yW3JZqm3rxhuOW9mFlD6nUBqg3
1jbi1gP6cUlG8g8AKuJq3/fF70r4EpEqcQK4lBkt3HEAE70Sn/7MeEnZaSLJCwQN/T26ta8BM1KF
GDdUYExRwGmkhYLeFL2FaSW888kEVDi/mXjNYURAI75+oBizCuiGyCdME3gj3serQvkkRNhGGokb
h+VXZTYlRw4amxq2rVKQsil3ne85ilPWncGf1WrBi2+ETcOKTVf5E/qWsDKnJESUQHVEGMAU0E4j
l8wK7LQTL8hI7yqmENSwL8DsNZWQJ2gTfE/H5GuiToJFJEQKuaRYKPv4wvQBS2nBbAmFvpf46a0D
7n+t+8tJnsle+8fO9k/HgIlWJ4VeurUcGpH23Sw4s08YkZ1z9k/lgLbZrSIHodTysuQfMopA/mT/
cStesEF+dXhO/VffPax87ON6EGAL+88cn+MO4fFP60Q0Xs6PqyJDwizcSkEaxOKR7UIsHPezNZcv
x4V7CP3ruVdIQywpJqLhnx/r3HcYKXa8Tf1L3t8IERAQHTAVwGldnHroaUwpLtTj3alOGCHnn1SV
LtAy0vQgWQ+gmiaizekubN/qbQ9+QDlpl9vRrMR9NPHVi1q7SbDy2eW6ZYrndp/opu9iRaAVUz2w
jle9Y7uP1qkzDscWX8dxFbi6ZFogqs/JR8P0b2i7HbKigW8kRTkAyS6sNcqEvrQQSn+cA3stqadu
j5tCIi6jnl8f9WiU6MwzLSy6lp9BrJDZCnijrB00nDgXLzE0ZGo8coY6xA4g7ko05RdV9sAPbGg1
YpZhtdQIrDdxDrA5bTyPQYSH4gcs9i3O9KNtt2jedwbJ93HSQ+wifrpCj1JBUJleZ1KWTsa4us0A
X0Ecw1CX8MGcH3H5BuXLIEO1qvYqGhQOO05i598K3/KBPxSkgcp/nnKuPOotpNEjGhTT1dJ8659T
h1b0TL6djYKcOSrt5bIy1xt1MODaTivLy5dPfLDCikLTw9H+l2a8WeWQnNulR+Jk1Zc3nG9rM/A1
cTRWuYQYo3/uNAx0SHTxoSD/a+VPjEt9v0gxI5EOHq+eTP2sW97ci2E+bn9nGoSUVddj4e01HJ3j
YDfm9PPEQlJ4LrcIJ6iQLJgkZaHxamCABRLATb2csL5qz2YObhxA4FNWa6O5OgrpLa/9M1BKYfuh
8iPfElJPaw/ZaG6lZta2kj1OgzabPvvAaMeqPBSAZ+P+cS7uBuXJwLt93Mo1irUUsVDFmb3xfw44
Mv92qnWlUANa5k71Z3EfLDC+NjUvWTzYpriGOMlU+hh8lY+WQmSIfi+Jb3LR8ZIcw8ox4aiWSqfS
F2B2FU6hxrWMCXAuC8TKvM34fk/yDEm9LPxmObNUQGuhpF5aqdPsJ+57eD7pu0IMqnMoLkjOGS6B
j7DesZoJ2lsn/pG0jdXLSBzeVUGX2VqkWF7Ud5sHs/Wd31U294fnS1yxQqx+cwg+/Zyf2SobbClb
DVx3wvRbiFlE2h8vK2RrnmeYkSXcJwKFTyrB6wA0c7lVCVo237CCETLmxYN6jhT7k9FUSr2LPqoZ
w1xQMJFQDWPxfRNTKG0vesZmMhM5eCUABResBCwRDGHfe2wGmwluIxcTwmUlAFROfTXozEvLmgOL
gEe8Mbh6EvyztqJak6dpyhgePwpeqShqJXM+XUG2m420WFFuMCFWk+KrS5LrmNaSd23L/cTIyFWn
wuHOeuLt3WIAgB4zdDBdiv2kLLAhSs+y1SqdioyDvGbtsiQfeg/oqIzaoi6BbRqPHU6kzPsR+T+Q
rNUH5u5xYrFIifuhdUGi+M/pSISPlXIiNutwyjn7uPnXsN2PH8nr4cqvOtP5IVxAAkk4a1P4ot0c
n8+/NmdYZHhwCRLot4B6pocu+0HtmIBveSjUC8LZPxINt7IJpbfVC5iCScW+AcMiksXDVS03YCXl
4AD5ayeq1E8F0U9geCkwF2ssVBIOlduu2jHgMwOmGQUgXdl/iBiL8DVhThlrO+HgHNYzSM3CJPst
kEA552thNhqguQZ7pvr62PatlKN2t7yv8o48aPNz/Go5/am4OiJl4AD6Cf8+UN4W0ecMjpOiS3DQ
O3L66hObeNn6NQFlnmg1sFUp8Bit4THnRKOKZ1Rdq+pq2iKs4jqwUi+HY24Jyl8Vdy8rs8mEUwso
bV0ZAUATghZL5+ZsB4xhVzieLskYVRYS/AWQ1nZGSUljb0Y1XCroSDDQICyXLlRRuV/1Ux6CB5wc
5u7W6+ogQGwB4n29rDQ+aaoJ1a4Dl51TLuunWJHyq9Nl5RRUYoBpnziOc9XBbyB+tva8G9/ms9BW
FKpN5kxeO3IfC7YLZljzWmQT6NvCaGlvXzGC6ZLkw3PX73VZ6oRkx3Yn3otW8nVdpdtDhmmaaUiX
o3oEnIrpB+kXt+iC4sfV8tpbvhiwyxJv6/ccZnkj7T/61eWzEn8si3m6m8UFXts//phn/8Xq5kVB
jBvC9PZQeryVGepeSo3DFDgp5Y9iFPGTpOyhiIemnQRAIz/EnEAO0OxStCqml9sSQZkxcm9EvfTo
XtlsbO4JNdStbMcjo5Jdfeb3jZWUW0jScrZ3fzA89dmyce+vuz2V/c8V4hj1zs1lhuMGXvMaE+Jw
v43Wab7xc0M+6un1QvrZhDQMN0wpa9/nVXLtVCWOzX9XlQTW5tA97ybPYq4cc7Nn8qoEGVLo2KCe
xARX5+w/PfUCp5VyHiK//AAUg44mv6lVVNSSMeVZb+2anbmm9awiyaoWRUhzeib1Zpca8uCAte5e
mj1m67t0tXyh0zSXzLboyLFB1Cw/m9po8hJQMqqcpCbCAvFORNa5sbwVTfgoTrg1HhNfqFgQCXqN
lyQgl+3V9MCWTtkWrb0IBWoBSRa2pgw78jG8vT82nvAM9SRtgqbKyq4glDQEr83hqRa9e79gsPZH
FkvVB53Gyzt/maqicsiYozIW/fnmu/LAQZs0WTjCWzBieBM9yKub/CwyiQImr/JXsOzyPBRw3zdT
jGUmLW64zD0g4QugM7zo534y84vjEI4ZJHHXqSGl+m8g6QFdqgeeBThpa1jXfmPqYRoVLxlJb2DG
CSmsE3izRqi6H8c/Puo0aOUCly9Uvi2aqe1/rsu7ofYLwq1YRJ0OSza++0LCuYrmxflC0sTQ43j4
/FoFVYz13ixHr4CkIMDuOZe5BPSIZ1HVRo+qZ+ygZ80jWYhz2IlHVpUQYNKJp0Ljzrh3GvpgCWSD
EkXKVGwP1wOLl6jUGpDv7Be2DunzEK+EJ3uk5lN4DW+FlJ0JnJPzRW+QpfSupP3dGHng/VeXRfWv
7fEKOCYWwzE2E1igUQXTVNQthMf9YecLTPuQMWJfmQzQPCBFLe02KB/zCGrGpUYzg2ivGX9pyXDX
Lr51Z7oapHjUSOri8jJC9PsBluFMiYN3GpYv19GVd1X09aaUemefOF4bE7uOZqeD2pfj/t4wrh7O
O+RDs3kRfOM/XfY1ViOFSYJZysJdRR/LBEUTk8r0GW+qpOEI6bfqpylRq4u8DIg8BkMro07y8r1+
yCgFq4GEYayQbHx2x9RHF3roOhgHAducyclQZ7Uc5xqpb+KxY3ZzXw8seXv80WIymTiYXXj4dhS8
+S75XXN8GYYKs8lPsswfIGgkjMy8JkjdjqmEl6I6Tp5PcPLWUOalNH7+5YaUmNYJZdo9tN7vV788
UsvQcPz/+AvrHsmL6Dkd3gip8y1PivHjgi7KmZ48uR7XVhvdSZ2GezJbZzwUDieFlTISDQNDQMYP
n2VgSpO/vBC9T/ecEN5m739ubk7fYeRzcDHAl565BWZT0x06xvQ51XKvyjPe7hgMItpaC9JRCznd
xrAcWsk6GkEw7T/ozIWxsdsf34TMxTczr7q1YkpUIkrA7lP/ew3WvESnz6bbyR7k8bvtKod7B+uM
YGhspZCWBqd3bEGc9famS/2PHMMu3/z7+p0LmcVn/AEcYUjOJxnJjgilwG/u9XSC1Isd3da1/O/g
TbyytgRCT7bMwL3i5WrWEHYwMsv9bjF6fHtCVc/41FcRWlNDQVb1gMr8w7GNhpVkmC3JMd0g5AJT
nUfppQR6HRBxQtd5dIebJWuGXH6F6BgVkhfe+bMP49c4Tziz0UcVKhxmYuUO763I0OQ17KJV5xtY
p3fW+/+gsO1X6C1zUrIguZ7jOrRuC6c3zrJOtuUdjaT9Zi+jqQCeKdaofAaVLeL+OQ9LqX7w7IFm
AWPuC6XO2jKdnIPXJX1WiZJuVv9mnov3x7ary7VJqyKJY7s6UGlS7F1Yxfz4rpZUGe4LHCEwFFza
UeV1ECUWa4hsYuksr/54rGA4tJJ5mH8+EDh82Er8aVOb9Q62YZBS4VjuuZpYLZtHxbzoxqn7cXJr
PJNClzEfj8w2KtG3yuGUAUsG4wJMds94++j2tmil6iFWhn0kemYcASKTcBpjDLEGm+AT6/PRB6zb
8Vq1cxgHG+oieP3j5UD20J/qseKJv0erd8W4bvXqKhcumu0f9P/6qcAly0VCQVWfhJC0rn5aGk+X
AaU2LkuKuANnQ6klLaaPOqC3SXGHvSmWObqNcsTSWnYVQCsCNfiT9ORAhxQtLOgiAyn/Csz5By2f
vPX5jDrcOyKq+ODEe+u8uYzBtgfR8/gvDf1CE4lORwqAlRBUp8uIitI76TJUARQR30Paspq6lwd7
pSXRh2jlZEXjbtXmgKzFGDsuxnEEfw+pnTjJ97rCsrV7Mu+bpn9qE3OCqvsEwBvvYegrypexKBm2
513zU0Jlxx1ZP9rFlg9ktk42YvcQGTcFNjixtX3dZsIuget/PEQoG1lwTCdEiid6o7g30HueVfU3
pouwx8elOaPX5pKZF9bHc5Pl6KW7uANWFmh84fe8E42qOilAHACbrNp0JmXPrMZ0QSoTOokGxWx4
SPbBnjQB8mqY+VVZ407rWGS6yjOryk32427gApbPjCvZDdLfVdo5KCNC1PSpSK7wMA1WSNKKN5q/
m5WTSbD/RoMvNLFXpH3Jb9GY1WJOKTQCTjo4M4T2MWY4ghZrWkhJwVieZhQYJctfGg+kEQBv8Dfi
7OgagQB8E2KeW/x/0gd8C43hZwgcSKzng9QGaCYnnz45OWK0Qh2CAlJ1p4r5ETsrtQ0WkijtTrZI
1H9C+RskympMVsfbSgLvZ2E0XewZCZQMUQV4F6FcJvDLTsLuGEhTvqqJLD7JC3maZz0aUXFmDb0l
qx70p0eTQBYeK/qWV1ppF+c4zbAZETpccNqdFA0+Nk/29l55oYDmXvKIq3w8kla56dIRoxK5HDbi
EJoxD0dzl5WjKmrdzJUzWAtM6p6JYnmESNWHpFEVWZ9dkPEpecLlzbhOupagLv9wJ5OzuKRo1Z+7
z3WewNfpvbfx5maWQMfCTOV/2tD3mE0rWBGZpLqz8JiyoRWonV9obqfvASAVFBEJ070S7pVfOL3q
ED76L0vFe2zM5SXHg352bPC8TOXLISedQ1l6Sc6A6eluOj3SoGj5eyl35fxvPkZGku8fNy8dlJ9H
MB0Sy0rX+U4TPq0jz4YnI8FOrZJ1g1qDQKTuaoN7qBsqcYmTelzX7bMiD6NrQmGh/2CJiAUrjoq2
ElsNLc1GATC77DBP4FKta4NgHJCIPFgIrtpejQWGWSF6M+wUrS4LKNz86bMO05R6m0Xp4rVfP4NM
wsAH5Yf9RApvT1wQ4qtjw94RCcBV1Jltzolad62OuA6b41soLp39CwHNJFqOj66DWYZzVw6+ROdh
bixaAgr65iXv0DEguFo57Q/GfI2JPIKexjPDKL5k9/KF0II5HLFDAMs6du8wo6YWsAQ9gzAoU1+J
aBtFbZCIId5Yrt20fKbLwCSVZ3a2w+VBgSuFVDPL6GaZJCeZLCrZp4F1H1Khi3ishkxzzt6GOSNV
eIKp9taWFgCCQPqARdbSEWP4glWclYgw380BYNqIE8i//3O9eXACQRK+SJy65ZkVcQ9At4vfti/P
jjYRymxBgkaQqDf+n38fW0Kjnz98PaFNW2YvyknQ9cupjCDUsORJ+NLUPVOrvcqslreCjRcAPFXQ
GwjAcnRMK2s1Rlp8H4TB9ItLutOuKrsqY7ODMXQqd7Svf6UKkSkOwworpZwY2hZn5odRS5ZCvmx0
KjqfqFAsuXzmnLpgXXe9ieW9koMl/LFE2o/hrtT491mu23NBOUovDfEf0gyfLRn9Qlp1F8dtjWRT
VYdtmUDPMeu2eBXTSUkmk0LYlsgLKH9OyRQ//IW+R5dWSQDCo+MMgwpXAvbNMR6KJuKqU8z46RXe
yfC/Jr4R27tvhg1qcS9WqGMHSOeX6VM9c1DDgVI/b/UxaN3gp+XxKWhe4GELyj5DNcxHuqUTjcLH
8WzebkPSg5KEYACQQ3VHm/SfQKIRyhB9N/dXPPwIv3CnV63wUN+NZsLmxH5+6H2cNGUe9wET0Vt8
rdKE/ZYBAWwQrACFF/uJdd5IVLd0yCVNqDeZAD0GuNw3kOB4korj5/N+lhYMBQ7NytPrpGR7G1ep
ks0Z9qMktc45574jUn6XACJIfPAhUK3TWwDan2st2/2sDCmNrjz12VGH29fx8BnAD4FUJ9YlQp8a
B+guM6TXiJ8YffdTing5Bc6rHwwFvpK8Ybx5oDpWLNM28z7YEAmEgsJUivXhlswL/yjme/x8fE2A
GpWj39fEXtJCrStNkQcBLhbcOzrvkP6hyeKbc/CSi7RMGrTxdGGSNk+Zgc+kjM3gWRO3Qlaxgz9W
f51TyiUogEWViXxisqAhS91vmu6ScbVFsuhRihhEUNQvogh8LKsXlD2h8OmYbfyd70hvWTRjOg4v
2iApwdbtG7e1lNYFJ9Loc5+2YJylZf0mFUHB8ebyIV2PDFJR+/bsd8Ep+kuR6DzCJDW1nOGKqoAG
2TzVKU7ASIlnfPxor6jRyvMI/O5nJxutbqIkRn3xswSAVa3V6fKUkwlfy2JwTYbwGcKIXZu0tMAp
rq5E6ndYwkPbmcCKwVfpm3vkAV/RKTE3g5TPerGcZrROBY9qQkKGSjvhUWEtxNrWTFvbCfD1Py0a
XaCiz5ufJuuHa3nZvDeVw8+yatbZfagLQnJAT8IewtftdM5Pqf6fcuOoDnfuqdWnAbqf/ciRfWbt
mVcaJ923lvC3tJyZKLDhT9AZk7txMqVovCeX9WrKgr2R/6GZuNoxptsSXDMmBTo9lNb++9nehN1N
sRlXaIvIORHxVLw3YtXJ9fdgTZGB1+EpaZD4rHvEGoZubngL33uhClTJuWe4UibnSA/9qONH4TMG
KeAZbYRV91LmgTXQ9Ys/jDaUXqXR9qgKMJWzWNV57aKiAHHoGc6zgquQwFoaYxjFjr2FyVveQeDm
WGCXQgbrFenCBPRbenOziaYd2KTm3sYC/jsowKXR8qvvFDqLdQNmqyvG+lSkU7iaFUZdPxxkoYsJ
JlQeD/heQZbgAtnCYCkCjS7P3CIBBnjeVmoDnq/Pj/Jt77B995bt//Kg3Qid3ZXg2Z7GC7DjuwJk
3Wc/4KPq+FgrrZFfpQGAMyqssIpwUxB+yIBdMw0J66S99xCZuHYDNWyk9tp+U9ts1Dluqv4u3V31
CnDLEDGZ48m+CpXI7+8Suo05mvt4pw7SpLM34tIfC6Al0nLhPrCQLvGCRoR4cTnxajgDy9NICjQu
UFH5T+5ls2PVHfbB8SNDp/+RuP3Jz9C1AH+U6V7uqB17DU21e2HRcJxPDUaBtqaMVXOGhYAdqbi4
Bxb+Qr8wdmfQ07KvHa2x347f6MuM/M0/nBSv1+Nb0WaIop94OXSl/o8N4JT+hhT3jTDortGfPTeG
i1ib3WiNhHDSIFoVfxurtW39TtNPNYdcH23bKwGBxms9W0N/AKdyH2WnrrNPAg8SRBgQCoy+uhKQ
3QIYIhTCDJE15A8ziTV+mCHjyu5hQSd2Whk/Pnx3COrfLRW1BNsEoD64DQLI9MdCaFbi6jkd02Hx
S1dpIRHLUnE6iSm1OQF5YCGAA3i1g4TlPjtb6umL0EOVQKMnVTdTLVxqrUwvwQ3PpYZHLXdLf8zU
/EPW76D+JgU0VSp3BokzjB+0dOWE8tZNZy5SZJ707GJSzLhsFV7o6IQE8+36vukP+kIQ/a4TmZBR
ooPopPqQUKaotCwL3F2YE17ZRWcl7qowzFIEcgDlLM9a/kPjsMmiq5vH8cbYsnnQSZO8X43Hbzu5
LBVg3ZwdSRDNCp8PAV2ZrTQQUIxdQBm+ywLYcA7/F4UqlvJxfEMY/lCbZ53/RdHl//QrZRhejfJv
tfSxNlEt+q4rZRLxAhkElRee0haOOPCJtwPIcY5HXNOofI5UzJnS788QNJLlYYuZwze8ErH6gSZn
eaE6BbqdEA+aY/T8i1wpSjNhpuAHVxlQuBoYFJOxdFvRnYyrvIYIFiWIHUbKFMBkSm5KicRp6UD6
yHl9AmmKhmroNT5w4P8NNP7o0hLE//X+F6wXxPfXhB+rH4W1gSNtcfVrdIAhdAQgxb9dpSYKTzfd
S976PCvxaxy+j8cdaOx5pbUg9WC2ugnYnT7nIrdpZl/sJsgBEVdTb7tINItaEuUMVHVQ3bSXggwB
xTsV6Lj9+yJ8RCf8XFcQzHfSeFmC00YrNyxzEnaP/G6HxS9hQZA16fdvntj1x2lS5+GHlojSQns6
9v02z7PuFozhyRuaPVkBqmtWlYQYxaaVDAeewut7zL0NhOvye5eOtSq3tP2otO7+oS39ZvMefLyY
/TZba9bX0UdivmxgZnfE/cEijkCsCjNZ6ppclEBXBPqdQwo1YRsTCmhaFk2OSzYpT+0rdkU/Hmgv
N8tzCRjd6G1rKD+N/b/+90Z4XIvRFzAhcfoX5aT3mlKE+EJSsIq6T71kHAPvwPdMhvOtwkNaXoi/
DKiTspmq/nB2vWdVX4D/7HucCGWgPQ0xxsX94qY1/OaIoDHmqHb3gvBtuIRsSA8MEdbrfRIqbiS+
UHLr7mnFTkkZQncfsNu3sShKuoej5TrfBEM7funB7xgnyi+dn5az2knQV025hNflN9t1phDn18Pa
bGwUP8sHdGnroZ3y0WhPWp+XTu79vYEBi1pHcB3yCZz86qbjxveqNxXDP8Bfdt47TPdiS7b34ZO9
ZV+oipvdWCDfGjLS5vtpf7P4fuP6ML+WxSnRQPxvqzlpEKW355+Z/4aCIPFeZjYoGoaHK4WMYPM4
REHCRvsOEV7Vl83O/a8QVC6hbKmXI0g7kGV1HbWzFc7qNsGdari3VTB4eUAphir3TI6JOoxYE4SZ
kGFJO7iIY8mRsyJhqG4UMw7M8XMp9DNS0j8Ys2zdPfHyJD3Iq2Ycp+z28d4OIgNZ5Qse3XzAXySs
6FH7MJglBB6yLbWXrl/lhllwr61PBR3ZXfL26FsO3hz2ZRWrbbKVHbcf0FhFh1E8MeAaDTeiXWj5
ZH4a2c/2kdLX3LoHaXNqHY0NygZN93TYct8TbI1+PciDdEKI1kI3La2g4n7gjvuszu8DP2pAktCo
EolV7vzEtyK6YW4XM07/cpFuNNrV4RZkWBd24FNkLPWTxw1UzS595vBqzIVtWlr+3d79mcqi+tC5
xgfBFXB0en9NO3Aavxs8U+OJhNVSb74HUnRGwh/giU/FDyMqTdacyXk4O8UIDxC/xD6UBTTbzlxw
fsG2H43B2r5591c1H/QRphcJ8xdqIy+8KxDmiz4Sjj0I6fsSrxJfsdAy4F/QmL5H8E8feQp2V290
Kjhwhs7lEVBppBtDtgYKytEq9cw/ADyN3v/L2r87kTPET5Ppz/R60VHtJtCQirzUVRIhqDpBpiTo
ZP6ytBQ6VWbAOnYMqw9pkJXfvSdtvAYScEX/lqpIUZd+Mi7D4nTxX4bm/NOJa2oBnzwRuHomL7mq
MA+c7kQLwH0IYn6FzZ22/vHJBDICfky550zvbRdcfle9Jl/uj+Mlspovnfm7P+v+P+5nOsYZo0qJ
hn80MYSHZWyfQRUpbo3SRdkQ5nGq8uhiSz1LQL83djIIqxV+2YmuweFD/3a+rVkxe1X3+UGbtcHJ
yOls/T/xPCA2Vi8+4VClwov1OF/qUB4nhBt0UF/Uy8yvbw9v2VmGc8vIaCni3uMx/Cv2vziCh5xR
W7fYSXCH9MPh9K8zyxnx0rZtMUNaVqCpzfNd/qnHO2CezOOhlry0DPwX46+vc3mJXR1hO/5NfNgR
Ogku9xvBHSiRKoK7ZtXyByewG1aq5S83e9U6evx0yw+ChwOUeA4oPq9/ZCTJkamUVKSYL65O8Bg3
8NnTj0fp0g68GMlidtCvDfNouyNdg1pSO7DEwbXDniulRwXn3q+vthFV2H3AMqaah8UFZsii71Ub
S3K3tR0oGFmjju6m4K6G+/qKKhttrqP/AelDLWIrDb8/76sP1j4q3speJaaiYl1ERWkp8944hSiO
XSNX31i7Qd7EE/PXeAS6RdjfAOf8xZMsKzUPufunvdaYqR28pBrUUVZJwN41QhcKmV7eIDww4Iwq
BeZC1s3Lu/OymMhGcs9VKWCxkDogWKUwr4kBzFwXDGPjxJpkhzpcrlpD80gv0wcTJxGJL7/ZOHOa
9LaIzGv4cXuxegIEZQAYZb7ooThwbv8Aiwm+HA2gxI+fDa4Fcxv54DE8U/8A2G/cMpEc+Vt/w1un
w6zrG59YgXjunLf7vfoHEXeZ8Eqy2I/CnClI/2Rbk3VcOkaLC2Q11sWCmDo6D/tl9mWs34JDvx0C
WCQIeZVSDZ6FtIZrusvYyykFLPNpVlX4v8amUL3vgScv5ezpXkyZuDNkdFoRvvntJQzjApqxN6ha
C77TkrwXe7kh71dm6qDPwDHWPRW3UfjfmpBXS2Wwh3viB21OoUpMPfsv4kg/G0Tg/ec+om8pPIJl
1WLVxc23FGtK5zt75iYJABD1D+SYBLJo2CT8D5t899UZj7oQCycH4qHtS8fzqC3xBLZ2SplO94mA
rKMDTIx9D7SFnBb1W1g5Rp6yaLp3lMcSypelOvjtX7TK60jTD5B7tvnyth27x8hV7lgWlg0++/bZ
My/wOev/vASeJBV5Yo3VE+gI7b3CdcLQu3HZoKuYo92yrPKsflcA+8kwi8l4Ust14wzGULCt2hkH
+V418/DhZFIFdMbjChI0q8i3gVYQq5gX+vfyustyqIiHdK0eflxqRqftakrviSODnt07hCliNhHj
+znuZNMLBTK8cA0dkPk87wH83kRF7puUIuCNDtXELj1JMr2UEi1Mbbj1Id6DQWJQnZFLEy7Hmi5T
BFML/APWkmzPHRynx8Qmsw19ymm/Up3KQFu07fXUmHUzPjSTARn/AA90Xb9TPoXJRPTxqMVuLVb3
DIlxWHEfHZHAr9AZ1SADjnXiX2/S4mTOaU2BzHnReEqMh5eO9jClqA6sSMyi9VO6bJlTqHIDdHCY
GAeLiQi5jEBVmr+hFAyhyEiukczIbo6HcC4TbM6NcgYYOOiYZWADnPa4UZso5wWPdp+IMCFGiWLc
KPvlcZNkX4r4BsYVSYd02yOg2IqXJ02OERE9YZenwyWmIoAhybsJffal77KBlFL2+l26fR632EhP
Vb6sORTe8WQLfYrx3kfz+FOGwku/SZIv8s9F8SVMjiJtQ5nB1KF+2zARr8R3yLoZ2j36FxWkPiLL
HEaUx86yjz0Dku+ehY6caelRK8ePEOTvHNZn3JoLLBMTA/NQuwd1HtwSXpllHMZONi4wONCGy6zr
1KqOFvfuJnqN+GUsz6chqoC4KKSUql9llWQxO/bdHr15nPV3Sx9hwPGXa6XD9gOrnqiaOiX7Mgna
OElBgDsewatD6zCNmgG6NOrD5koF+UofUDXomo1sYiXE1D7nFPpxW4l+7RAvGQPRyg/aOG1JSpVx
r6lnaJTS3Vadk1K3B9bvU5YkfF5KY0/BPzGOiIDTfXTq4nxR+EIpncTP0ZXzNqqqWseJpC6kJyt9
lV0HRe5EzKcIHEmBm1lNj74/+fD7waPr+TyvoyJHOn69lTyJlzjz6/9pmMorf7cE8sORqMC20a1N
ZQ3sKdMkCxkuLbxh1Pu07Nu4dMf6ucQGHL4bZWMFJGD/sObj2AJmbV8edEPcu+of6Q5Oi4popGF3
Tqm4dpdgIrxR1QbIym/qrELEf8/PfyAALYyqrjW9LYsTASA4xlKFkL3Ewdgk4jyxkSCtEvwUVfqg
6WNGfCdESHSfx5ACX1cAjV4XfhWzlxMJBIMBNd3osr2tdsLLW7eRXotkYSpg2grP56rEv11Rvhvb
Mpeo8/KnYrEiLXRouj/jB0Dgcm4s3epNg6F+Fu9JidRnzHKInyW8W77ik2nA+ZwPCgIqNbU6IU+5
J4tJXK7XLjquiAZhLONfN/EzBnBHaBR1PKGQ5CMuKLza6X/BrMhzPmo8mEcZGJymGynmwpVEpdWo
D45M1tY+D5lg5c0y5bnfWKsrHqmPuxknngnsevxIOtN/G8ZZ2Ar3j2DF4BgSyopvu1od21zJlEXA
YcnJoDZrNUNYpMaTQqwE1lHFFwl+AjXsqJSMtNC8Y1ODmV+IYcA9BIUOjdIM/Z/cC4H6z9vUFVsl
6Fy64+Rsi+ZY+q/T8jtzURuyvk4VFu/dUMLJ1QPzK8YzalUSeMXI/Na+TVJJZnHKPJ5tL3VX2CpQ
kuhntUCd5xd3o9F8+2UxvqgoPffqhY1ZbACnJ5dlGIPpIzZzP2iz8u8Nkt7o9b/kvc42Tt/R2lL1
GRnpNi/RRp4dmZG0OsFPkLJTYSWIwqmglQYVURQhRnMF34uqQZUVePXcki/dCFWer48vkKKx8xAC
Q2MQa0/j9LM2cUR/zpLqX3d93zmmz2Y847C0yXNObOmSChbvKCrfnADiEwQah/zFj6v1bMyHdWo7
zwvCiA/02msga0gatL5JzrGzL+dzGzSoi4hHFvPUi0RfAw91dmpyX4A92SdmdSmCwwmihZOIoi6Q
XBaBNTuCkX40iejbduYyEBGvTxUWCEwHlgq2974OLuRMWA58DObcLegfqGySXGinQdTgXGdVHCil
sL0ZIkEZbCbDhaclHrhAWh5EeqvuEXLzjOYp6aiSARAa7yUr80lerN+fp27Db8GHQeWM4tXMJWxF
rp3Y9/CaMFrVpKDMtyWfylpLa3Gcbskwhuk8w3q5dTcDzzkjRZvR0X8H4JpbnZg5J1abjutYil1e
bN0Y+WqVrPmyeDQmHThVZBvx0D4QWgTXMwUx7+hjYAUT/NTh3tTYwpe2D30kAgmH3WOEmhO76BA2
ROq6qI5VX0gRgcVdil5YEdIXXh63inzP7gpjHaBqTpnWtGEJATF0NXTH0HDIw75eDdBr+yugyxSS
Sng+JafLbpzfbw7CuhMccUB5I+fAa3F2Uo6abWQhSTx9ZBEeBZ/IejLdsZVRKvL1MCk1FNyEVHG/
CQvy9QOGLpNPlDKJT5f/xtmoYhPDdIB+uyU/3/L07GMEmcYskZkR9TYcC973qgef0/R8gjg4nQur
ZOHb0/k+JfPdM9KfilgqJEfWrBXQ4Zt6c62KWGsDW5Y5UDL7ODwlS/hPFbyVQSL9P2RbdgOeCe5b
klSof2JqYtkT9t6eVL7buDS5loJKQ02+16XNINK/y+2vNoD5nDRnx89U9una6IuvIaejlA+5s2A1
3A7ETS/wuRi1LrwhiDIn96D+2YzY59lKshH8m7htnOfeeejfIos3+QSxXdaHzHZCFBqfbMeTaGrS
hGUOee8jIG5P3Wl5na21JWuKtbMUPuvs8zAM7WInT1eBrqmEf0XEJ7fJGt/zFcGtsnNU0x2lhH1f
vVR9GXoqro0gcRS2uW6dxoNBdwwZtFYEn+m1DqCev0bLSuQo401Jl0RoCsi/3HNF5xmy5RzkOk4x
Ub5YZB6MOww+CkmHcwtFK+8DiYz4WL+yLdIwm74WK5+3KaEilPDWR9irNje5HOGzybJcTZY60jbO
ET5Y0pznsRTpJa8v5v83jk5Khhr3OEzoKjBNVWPf4g21sB8Z17h4MtyPUk4fDZZjsmWrFiuAWEn8
IBasGd8IobN5c0b/H6FX5QK4Na94c8mIErH35ND+fRYo9jb7ImUBO2QBZy5Iv1O0R/EgOBKAna4I
U0Jt6DPFQjB+qMkG82Mn4EuuYIln1mq/uu7DGLlMrmZHMvnyBCeHIWiABBaf4WfCDpf9XTPpMPd0
oNv89CG6sBqkv+EnSWam5BlpjL6D/xsKFbRtevxKIlkLa45WdXd3Q7HOoyOMwz0tRB7NNiP8Lf/8
Bwl9jV4iZvedGOMCcWY5TZDcmve2mKeaYL//pYv/NtF9xhEJkQkYLMxsj6tUZjYyP3VnQKVZ2oUP
fd9PvROnjHiJWHLrDXhuMZyitqxiznn2O7hB2yEdnNR1xLM7kgH4WdxfimuvMpKWxwj7ineLNEyd
9JD8/xawtdN9YiNu6OuuaON3+nBDU0BlugpD1FJZ/VeaHJAHi7Qpe6CybxixvW7EhKchPOsYDqgr
T7Pv8su1BA3vPlUNv7Hb5v3y7Z0v9DjJR/kgAgcfJq80Jq7pDU06kJ+MmAVgYaq6fjXImwQih9DS
0CDkfjAdOUfVMFw+dMS9I4ALkClMlgHBXmVXVpwWq7QbHt8lDPC35CJWTyll+Vao9Rqmup2/qCMn
pitHIRqKx5aE9qxPMiK6zDSl5u4JDuTva+1DFea/Yaqo9eNEG5t8p478wDDbmm+HatEfcZqbQkj8
58GxZBSmcsyuPhxCy28VyFdtaIE1c0dFL4Q+phO+AJIFYUsyWgaoA9qA/zaSj0N5MR43aym0bu9e
351PYbmocZy9/zEGNfU7pv63mgviTrckRBHXi6fdPenBeMm9UxBRmqEWETouddadrPJT9IODi+eG
uaJxbREyirGG6812Q1O/CUXmSwo/0fV70xNClvuY8lvWD0tA7IoDJ4u5b0FQunlb7OIK7ffhA4lp
Mkz4nz8G/Xx3G8WBrmhkTGpxzLGH2UUF6YCKip6pDUZ2l9M8r87D3HlJWOpV6EStJXyp6riR5lGa
H1d1JpT+pYXcuER8LBgukKvELC5k6PUsYRbvqHWnKtAu3lqaYDxArQ9O2ygC0RH6X2FYSxlzVGFq
Dbf5ac/pUtwXFXx9FDQisHt95Zt1oMPB538L3K8RCEm0qXNLzuNUVzQZyzIo0f7XCJOzHEHFyP8h
2dZ9eG5WW31YrESVaWvbGJBOcUBHPpUhuRS1jKMGxca0ImCanYJhy75yHjMKJyIMevUm5Ius3ATR
7SlgGtCpxAF04xUOPddLwb2RKNln76t7YaJZc9nkt9TRkhMNj4fQcsgSSmwTwYBpEm6bxDX8wUeF
/HgTNR9aQD/GQbv4DOpr/dSxjeZ2rZURN8e/3W8bmO0zyLrnEAbh84U0pL3EEaATt8Lsaf8FUOMh
sqX/A9u3rKAvtqcu6MmXQbIbWZL2n9eaFaK0uW6itRk0Jrho8TodyrrUHqpEq1wHLsTPIUfsGS4K
Od9au76UYZtqLN5j/qmRd+rn4rvsRAsNPg8o+8zGfMVX1zyoodcFXzTaHJYSGPHiYias5Rv8nfuj
I5STfei6XeL50SPpaPFeZImYxT7q7fq3ORx/KmeOOdm6dvV5Y6w7seDt4rU7KtdpZh2GPPP3+b6j
b+1b5H+FHq3PDCByX4yYsgzGIFs/pvRyApJT3k752JPt4e7+fO+LqF05crEmFfrpQd9E2nDPOqNo
ughQ+ahiJAFTc6v0bo59Km7JHayN4zkTnMOA11UreLwIRTBW9DmYUkBQ1EdeAlURYCjC2XsDbBIl
B7s0YaQjac4vU88DBv37u/pqVP2nXBuDnpqOFdtGwYRdxb4y3RqoQbIr5KKxaFGM3Abs0knAEI+Y
b6XKPfssuwvh+k+jKO8IWvi3d0mlBFG66QSqqWkmBWV1xuo1TFluA+HAQbYd+dIZ96b+zISkySd1
G5f4FuzU9xTMqEtuB0dFbqhilGISKJWBXAzZJhGlKfAvhrRHDQ6ofwzMPAGR1cjY2N4D71P7kymm
uQBgqWybkkXAfMe3d+f7LcJ1s++uzFKXFjfmBP74IfLxQHP3B/cFOPTJJCeH+D0flV8tZw0sAjTE
aSAzOhiqmUXuD5ccERdCxAR4B8vrB2pKRDpzSpyRjx7FZWy0XeLtt02OwFPKHm/LyDNFw+QAX2TM
TAhlf7cpjMWZXTqBz/0ym3OrgIuhJldtnnh+b0ap57JdMgQeRnu+II5PXWTSqKpXREeTdmz39ZFX
WyfFij/g5xrNZStmkpc/YGuPuL9T135Gr9PwPxxycAjnZZsIfMuQe9dRoX5zErRP/rvCTlIC9GOo
qVG/rUDkTa0GImiQnXZzJic0AubxGsArILNKRnr7vjUvSIqaQACNCZ49Rnr2yioKnYwp+GjYzewT
NK8Zlh4E34e2J8j9LHTZMVLCigC8dp9eCY8WpI5u1SLss1yz37vW8C6/XPbxAkG7SUoy/AQ4FKNy
c88VJgkONgtH/c1GMxmwMgOm/CG8/DhW9neqCrulokiyuPJSaY7b03ePtUITOD1c+uRcQ/soXSv/
X4VNL40OfyOpbzzFmmuplXYcg3jtcvnXcDkcz4wei9SkNzGhVjbNtucC7AwjVwk6Nz8hUDMOIQq9
5gcinTG87VYQ4N2zFMHCii0uwoMuTRCXSDvylckWYB3awfLNTigsBO4VmCbGyAZdrEMepB9FhLlY
ytbG4QLdeXXbf01AB6WaIG/jrWaXfVU00PdlWcSrIDtrSxEwQiGRFgTVhNMQ3madbmZ0Uwp3my3z
fmf9ldfBnzDsYp0zH+posSjNsYjd8T4+3HVTYzEGi/H1p8iqfHS3yctFnn/wt/PgJSFvp14z1xVq
T/33ZUVTK6FQplcf71KGhkHIQDe32N68FME/dOVZVDDyvfoC8r0y/f4IaZocifXDvGnwnf/AQ3RZ
7eBgRn94nyi+JTOsjYbY6XR7eK7e5PMSrNUz7CiY6Xbfdv6pQugHIBqAxU5B27o59ftz9BQ0/T5a
hPDSODrKaDAFo5hzpduLMU5ajtIORxvHPNTsT4qGUk2iSt/6hVZURUo2k/Gj1NQ8wwKlo0/qnq4O
/CLYiYbK9/7BoRHquoUtkOhXiZ34efgq9pCDunLFXZjScvSdf9RrNHga8x35RHAezYHDrX1kO5xv
jIMnQNjA9XfOKuARhSvqw5r1EhmW9GWhm2nJcCC0gAQsqSMl412kafYSPzkvqecolspakzWHSNjS
+HsPTmvnyB5DqGn8L+QGY7MMDGTtB8CEplxSa92dNc/o3nwxvc3a3OPSekKRQ3XS3Kg70TPi/uFz
42Xd7+/7UeOGGkE7OpX/GKPrXB3HldWVLSVjJQ4O0Rq4pResFIW5cx9Jj7OgK6n1d+8H2cuLiytk
vHS97GEBELfXnUfiJiY08suMntA8UtQ2KKaN/illW7smd6qUHLp7mpHJ7ikBb05TwDL2UDBpAm9i
jAZEnPgzky1sRJbFkufsY8CJlvLTc2YkqjIE10trbzxhwvVRTxOyvClmnJWWunHLshfZbpMqTDhL
4ShJqjjD+IAaDOwbUv2pzEOrOR/YQzDKL1k48p1kWjAdzXwOMVE8geH4GsoipXqZcCwBMAzLb/bO
TBgx1V+gQkIwoLxI8SpRERMpAAtruf1Tn3VJndP6/vzr27GBHgMHlWBVSk+hJmK2IWH2bSYfC1v7
MwG3nCwZD4zkGKiYD80ss9ys1rwmLRCuPpzDNqcQQGTxObQ1wBIkUgSIMfMSQYMqsx1GC2SjC47L
R6iQLZ97ZRa9RQhGAwzt7nhuAaLbvHai4zfNcy/Bj2b9WVmK2IDzpV+D4bU07/fI6bIxs5Ef35xA
6T9DYDsT4iSJzuto28w1wjNPQlP2Z+mIT2VEZ/6bM9mFdMFEuhkU1tVus4Ha6i/bAfImmgSsX0Vi
hBHgkTjZRyB+zdB9LFcktlbvVBnmzQTgMQCxzlKU78uTLhztEuWxdIXV2BK+nSV5ygIXWUMWSCIV
7TOJ89o7h3j67wEGCRY07SCA7OHp0mpHYLfQelrtYitE64TDTr5PKx05NEVgs/jc+QXgwDQU4eMq
sUyWUuPHUdlCOOY03sL20GUNLxOF07cRYanbu3Yycpdw2i2BbffJ7oCqe3srnYmQeIhVLQ0jgDPQ
J66q53oRYnCF+Q/CujyoRdJ+k20YybpLl+ge/M2mTFnnE88SUTuDbC7iJ5msdqDnkJZq12iNMorc
iJ5Ekdi2Es+IJNiJg3lVehsotasBRLm5KRcxPOC+BvMuVHN2p34d6H8CjpiBdEj3PN9ybPwHy+ho
BMMeSNdCN+DS+we6vC3WkwymQwmJ9n3V006tgDI3LbGoy2Ali3KKJHH5mTlD+GJQKmvI9nTvKHal
S5AWBSe1NOfy3btCooBlWtFlAtZh/J1Aa2oy4pzl0LLhZehNRFTGNi11g23YvMHo250wFKQZbIiw
hatmgE/lz2KEyrcbkpeB/nHHzGV6eUf2fpvbioE7buChaxEAPxoRpXp3tXHaec4Dc78KYxDzcrvS
YeTg3zyBBnyAkBfC4ldHY1h7/zv1/fBNKoEVU7XsYhz0f0YJqyKL8+TtWFX/9w1nI0ldvr/AilUO
Z7fBAQQMmQjA/ZjMdreCNFuEeHDegNiZbgRxpUL0doxofSkslNVY8wHXpt1Tr14x2eX8Ph21vCi1
fq/6dVX35zn0ruInYUnF7XG44/XQb4eJ5L3o51T3xjSexLWqGdk4VESlyGe1+37GyIg918/U3aro
l61THigrfIA4GlTbbLHnEK08fbTgYmahuexWFOafSmnien84KSHDPJBat821ZIlLX4IF/vTMN96b
eBau/aErtPQBRApIz3SUkb5gRSPFJtKS4GGIm8HBjQq+qDm6exU5aMaIb+iOksgtL8hTKDw8f6OC
5seLO9Q3409wKcxSR7bWiO5xizGL3zqgc+p7XhzALnd+O7vkmBwBwqDdoDrWzzZRN8GYqWiQP2Fy
DweVQOOuurXWBipB9pzCtMhp3NAkSra8m3cVCY6mEwXcEPoM3otxGzy0BYh4q6Jh4S2Fz/j3WacK
Zb78ivSY8n+kBBi9p3s6nashuP8b+83UOuoJOCO/bjuzehKgvaad792B3uQzO/8qSqIK9NAme2SQ
DL470e7u+EME3VY0JQy1Dh23Lbnq1paOXPSMNMXs4xZDtTa/TxTQMW45aIGn/jqIvhAihixhmb3z
8fuXiMPeJuf7akcbqY3HmgPT3sYFsKsYrrPDWW2U/LVaVwjZh0vy+jJNLFHAFBIRHOdxGxPSIFo7
u6PEMkFNsnkF50KRbCKGM2ebe8WcKxvg4as8LlyfpHv+mUCz2/D5lTPAeMX6OxNNbvEib2P7hi+c
z68LiXCFb+45wk71KcLepvRqrvA5s9uIGgLO8JaIJnTV6Ac/u4rZnbGkVRzABuTOEn7GIuTNGd6k
jD1EFO3TL16/BXxrhXdmlv3XMou/+M/nwzYeswIVlUQapQ6DYiurQzlEfXYHlajszLM6+RopL+0s
ZTfAxmI8MJAKFfDLIQdwNCchRE/JzjXbnRR+A3C2ZMUL+j8qArfpkwWHeK0wG3U85ynVZawiVVVZ
MgJV97x/um1DMtoqXNcb5+wKJDUVoYzYt4U/q5OPjV34kRVik+o/zcoExFr3Y6KZMnifPulVjvlW
c+6GUSzyDGZes7Drw2QVWvW96Afnqb/3ZNkThecmNRYlniHXUS9/TGYZCyY7BD2AS8p2Cnf+xPRX
JKqeenydh0RDlBYqpuZAWTifxPQMORJHaANx3vdJOkWfn2f2oxTMrEpQtKrBz+ueWfA8NdyaGCuG
iWk3sKHzAR8vqxQHm9I+2Y1+JN7cRq5fjs9Zaf8pz20yh1fx6L98tMgG+7p+efQJMO0mpEUIPjDE
xqUFhIrTv19gFnzP6N/qZ07XJHgg5WexstJBXaL7fjm7Hux9ZnKFcpSUQkya3EOcER+CPi7qXZxL
2avzrY7GSPPxQs1x6tz+NTbivQgKVhGkBrTCWQCE19N8CCP6E5k6VrObHBkP5voX+SfGowO3A9YQ
OMDjSSFu8KSSch2WzZIbOSNMv80RtufuKgxJKKloeW1bvEElQb1htGxm7yZcgpQxiCbp0Hlfk56x
SC7j0eA+HWFv9WgavRaCnuQi5X2z6uJNGzaDZScuGp8JpHkOuN0wq0e1nUPSarFfpV1jmqG/RCaK
fMnTOilYahs9elgXC4Q8T8S8l46/f0YsU+fjGhP5ciuXmzj/fbwuCZg1l0m7Yo0B+A5xWFeb/SKL
t9IwcgLc2LO5G8sSv0ti4gSOoDgm9jE38qjsbXcGAjhde8wYNWF73sQ+o3f6Siui3pInaR1Sqr/e
//2YAozEP7sS0eK7ZVIy4Ob9xsteym9eKdU38KPYZOrOnZcHZaoWz/WPMTlsWKHKeZGelrsJtc1e
S2K1dae+mKcnUQ9KzLnBwGQeohyflVOukS3eKHaQDETdqX+kf1l9rRVXcAD4oc5K0e8kOhQaWpdu
XQrbCdikN9Rj3A4xm/Lj4UnVNrYwnSiMCTm6+T+dfsa7p7o6nS+5lOILpA8Pu0LotXLXWRxZtE4d
SiTii3Xo1r+tnbkgJNbU7rQO0VRxs3GilhC+cG7ZVY0NpfGyWqZ25HUO4DwlTz8fNoKoghDFNYj2
d43gtQtk+/fIoOGoIB704J4VTfBMcD4DcLFefPbrRxxXK/mTtu+wdInPBbcBGFj3JxfAt/cySe/Y
vaga4g+YOvZE6xXifZw27KpM2jyrxb3TigF6spG3s99sTqvc7yuseIUv8VITnTIsgmW9UYo5bY8s
AyaN2MKSHiCP2yFgw023hXqfiOaGtMNtuCWpm7cdU3cmepSB2UKEPbBU62gpMU87EXbTQmfkKx4g
D2cnnTV2yJxThkBazHkstp8inwdEq8ELJTXLH9q5PpBT5l4H2qEPJs8kq9Zyjp86pBTTtJA7SIuv
QjiRXqC1CjWhmxHcGfYO6fTos2wMt0szQq9lWIWpLXvpIi498FtpLbzB8oqa9GWP4A+icxq9elvM
zfUZTCRW5TUouvNYzXSxZcL7I7Z2OIDRUVBgdcQqxDTeJ3GK56UxyqPyISFJnNbyZcGR3PAxYAFl
jEXt+8Lgg7CRPXWNCCRGqUb/349C6CZbeFVuDrCr0Q28QA5rvQwVc/COXF82DQFamo4sTYLsDD/0
awrwINxJtrJLl/hon3CGEluD0BlDS7zxrFbKAA/DVVP13fBNfA5zsyzi2cIDRAWjOTpBxer+WpF1
iBxQC1JyJFqAiREzHlhVJg1uS2/M+xOY6jEeCfEgTxrHMds1fJqQWQJzrTx/92YQXhS1tvvSv6pY
dsfqabi5dN6FktRzdAw2R32sAqvC+L6EIyi0uBnjOpWDs3nFg1x4Q6gvW+ZpzV3Hfn+ALkbfOYDd
gawVRd5gtJFNh43/xAvLt7nO52UZvuZgHG4Ifva1hPaRED8eT/o/hJ59OdCk1pnkpm4HmtwaXoLX
Nteddacbe/3yeP0ln25dXSskztDVg1R+TFLukccONv1/tz0/5xuiVaHKXUdqtE6HwxUTrooNd7i7
FjyvuTXB8nPyXQZB3qPKDoIwikH9QGHQFffUgLZdtuQ91EX5p53awn2LhFNcdNuMu5Evt5mvTna5
hCCx2ohlqcy3fJlGr2WkyPK2xqBraNboDVBqYM6JpMsKnajArenW7DY4b/sUNTyGc8pJyT4W2u4y
uGHLzGQEH7ZC5Jr0XiulXDD8fD+nmcmZkbFf+VMuqQ/e1Wgexqs2gb1zJfDlnQ49pFPQo+HjqG4m
LJBY1dGd2ETey+Nd3LrcAlYHjA5oCroRgP4VXV4opcp5GqlXqNM+xyVXHC7nLCsf9O1dOIqfR9jH
LbEFlIPaAxHiDzWG8hPUDoJQuRsMlRWw9fDQdKWJ/xaTy9pyD7oc+/Xxy1ZqtkAQ68xcAJxu+KXL
uAH6KIRgMcDulLMmpC1qRaBiyWoV1SlcyeMugz/0x2efSSXZmeQaeaFiAJ20Ep2L1ICE+/FybqYw
WeLA9VGAo31t/qYi6V/aHgnQii08nu7NaTCnPukMC68axpNY6/FovI//2u3WcLZpUWG17F6Xeb8w
HB9W/TmVaDyxGKPRzFPEx9kRpFsBnp3Wk8pNwtLKqxnOWCMtccbUIko2bu8JJKjyi5hoX9rrjxb6
AmJA7KYKX3qRmh/kqag8nx0PNilElLiicl0jdRaZ+NdcE6ZJWcVe2GT2EGiTjdbUrJvEunZk/shL
DutU9NjmzGwf9LOsgYxmZp1CA13L89muRqx0TmRnVddS+jC1xsXLZmGz3DmIeVOp3SfUuRZcHPI9
BpUFbEWsPO3IydeEOuq0uOa8kz1o/MADKAKWOIp0gxflv15px5kLGVvAjvT66S8WWudNTuDevwg5
bJg5gzmGyyitx741Q05/U076EKGrTcDRtt/PimkyWgnpCDXJyMJOH1vLfNvVojQ15tdNzMn6eclR
uc1Au+5qVXguhZw3FC1KA+FQRyq1pi9EwepkPH+UWLpfGzzltkLV6t7tgQGMC4kyV6u4v1LKyOHk
zlic7E8MNFrwbpfjfJ7Lvn9mu3Nwqp2OVQO4Rwhti8+TnsuXzRhk1uttxi+eQ9342oMCansWqh4z
ikBQINhVpxvgt/IBk6Olbh6WnLk7dWa7AG5j1Li6t11qcwkBok/qT1J13MP+ztHIlPEpR22g8USW
zKNvEeDBF08A9sMDYdTcZnpLbz2+ef83XieWj7aS4ON7GJRzV90SBhn7qKnmeJy0J78FT4n/NBEy
q6FjbppUg4FH4ihdBI2F0I0/iBa0R6//TzPGPUbZba6ws+JluPLZMCzyDrsjcisJdg6HpZHs4vlJ
p9hRB2BDX2z4ytzFF4RJqD/1+/twVUeMFJF3rAqGx9kVa7RY7bq/qiNERz1iXv3C29sUVPFEpKB5
+kGY/DzNaeS4nldnxzZlFew8uAWfapntB0rRjcqIqXfbur6ULb6U5qdIXv4l+S6JkIW26v5YxONT
SySefaTVxZ8nN23G9oIi4UlQB0bXzzfTw2sZowlyGVDKAD9xTFcS2mutB0n2T+gtvaIQlJ7+AYoc
ZW6YzDkL/n0tKupmcMatTIIzxar1rfPKPVmDJ2SJksO15ibCpxhqGjr+exGA4AiXQBAd4EUOaYpn
dBU2BZ9ZuwuAuoDRHyiW/JkkVqui68hFYEggScGUnpa2G2kJcGdWoSApH25GqFC38rBeP++I7ykJ
a3xPpxDppy++XXpAj3nPkoO7Xf8G1qayQHp/4oodEgp9hsotdT6+4GLnq1Ww3/rQ90Y8FAucAGki
gYB+NRw30+bnm3Ge09l5shZIWF1+oeH2Auv1grcKD2VF8tzFObH/Gi4u1MISMaET3Bbmpho1wD8Q
av66L7oV9aX3eR52Cb8EizJQ2YSQCuEMiWjZcqpuf2yqdhoHr/H1qPdSTh+Rlp651Tc/xcLmtDMo
33uXQmy0gOLUQtQwPMG0iKNq4GArYbFv/ek4yhfyQVbLioT4Kz93fcW+dEEWURE+yJUlam//ee4/
4BK/FsnftXK6QVC6+pIjOepb7IbW0aQDtkSqpyFv0O4SOnTbg06QvedMYg4IQKkFOd0v0b7VOqKx
mb3aSLNfFrC9LYc7fGnauPXGRdSCdHavuGsbu3XqqgTPYZFXVgh3/B3TrJgWNhyrmasO74SLbKQD
rhHTcbcglxjwf6Ed4m6HcKsggVGt6qkGOBKzrr/KfHqZ9ofrXWXmEVyqfVN9W9mph8pdR7WI+iQa
dZfzumBMUJfRYFiCJ8cxblbnUP7pDgIYTsyyVG0lxebX/HrckSkSibayQ7MobY/Gw6bsXDkGy1aM
qgfyXExgHYFWouv/CJZXsPs1Mv5vf+zPdDDSx1yB5/Onzex+i+CCCvDlrFQH7BzlGUtqEiOb3/VU
kJCBJ9c728OOaj8r23vt+4cJyQX6JoXBbPLCW1FziyBCc2H9a7XTFer1ksXJ3miwqGYS1/nrW7/x
WdjguLOQupEHBBicD/NTBVFTEThBxrib3+phzvWsb8PshKCHj/wa06+HMsGoYB+BJHsnYbcW7WTj
1t+3EUAR+cM48bcOu09+shbU8xuguCHg9KybRWSqyoxagaAJq8HSaHib9h5KkTHSwGno0vqtec02
6PCHDJ/KOhM4cVSZenG6adferWyUtEFlpFS77nqrsrWJpsiGYWm9Mkph4b1frZZ+5zbu7Zjiy/qU
n4Bux6dt4q0QfM9QDdPbNWIlPuJqy8/YsNH0jrzJmAP8KUXkCjny4LDBfoMzOg6aLhZhqlEGEqG9
SUogzNIdZVbf1FypWHlVCbMxGIvOjz+UnP2I4q6gkiFCPgxhJ9ZKPPsoiNC/sDIF/a7uPaEIKEzS
V1P0yUNT8Jz3IBLTeRpg7bOvKmxCW9A11c8gUnXhQqOEM7Qw4ujiuUpIpec6ZLtE9qA3ejeKR3aM
d6wD8OjN9uyi9XC6EQljKJZRMXw+v8xefRkYhZVTTgw8NYv+DZ+M9dlxGzcAfyGqtba1BluXTHbc
ONrW9m/SMwD/b1Ajewmdvz+wioasQpQIbj07+C/sT/THy0P/KJHcxLC50sbF+qOt5+xSxcyxrj2d
g7O8kk/oJpZBxe0r8NC0DzMShYObzSEAUa57UuJA8dClYt1DBWjPIhuNMGR7ya6Ff240A7r7AnL5
ZhOs2mTdB8SA0G+FT1YYBsJ5RY1KFMJJlNn4AOUnVYNN2Sa2mdGy7aksJfM3Jl3x1B3abYNvidgz
WsHKkhn1Pz+NPMgRffWLUfsnWyvAgPUyvZ00STL1xunkl1thT03qkILVBILzdH0tAOcbAymKM1Ho
aNlBnqQFvIe8sXHzjxktjMPFcrV2oN6c9FkfRku2VG3FrsG6oNZptO/6QyPfvvXITipsDlKNSyRF
TSYV1U2o34nPA3oPEzI9xPA2Vq3cS9jjBVp4VtLtx3jumfixObbr+ZPduMeL+aUJuQFi+vSj0nhR
VKUr/Wn8I02rggNpMAWuSmYF2JujcOzbzR7wdetr4YZyuE6dbHjP7ZVQbSp13n5o5Sc7n9ex5a1t
GWsFZGkcZj0vX7mPHxBXNE0AzOnTAZb1pqHfS7UI4ya+4F6vyycUCQsApmufxsI2C7mbzZBNUHOp
T17sUEoHJOPfJHKMJnxee+o4XxCUgN9I21VErcCwCm4eCB2XF4tCAIXMWHUwTC9GoMDHzeYyaK0w
tmmtALmHDbhHVdmMvx/KUUgG/TbgKY4U9P4ggEqCyKzGMqOM1WNpaPczDqIuPTEdv2WAsXUeMEOq
Av5GZv3HUHvUSL5Ty7OIYbUMk9sEkdArT64A9psCT2Nef4iwtKPLoVggefRwM+WSLf6OpQOYUV56
tabse/QN2PzvfDzHRRszJ5f+ncMzpe1/rvus99RIS0PfIJdYvavrZ2lAozrJQ81j2MqR7GZOzCJM
FrTl9QdWpLzlt79nnKgtWJXS5NZG+6t5LL6+eZxYSKmwtR2ppKioIDja50Iu9GaO80z7vsTscvtm
04TOsf6WSDvdBB7ggPeXi8SP1/oHHoPX7ircFLovKdkUs1jguQOSIEHwNfC5zGnADgIpPIU3CezB
chStVO3C2wqb9y7vM0SclNhL77Rd0K+/4R9miLW3mrNrZHAant/hp2RqfLzbveUlSqX4TaeS2ExW
9MWOPAAOXX1YVdwMQHDg4NekDW1EZaVO5gsAJOJws7/0SFIfZUN/ryxwM7u46tsp9oycQvyAYll6
aXXrSBuFxaq2V9ZNlUfZKkJHQgCzkoyIoPijXMKP0uZ+2/YXnW20F9PHLSslzFhKLq/+NOLxj0ml
O91ZLD5BB7MYG8p+0qkiePRwXrPbzhIl5hPM5noCzyMV/GTHe+L+dcv+NPU0pdhVHKjnv8zQA371
I0vJIC1lPPz67nvnpnbjNTraFRuSu2Y87k+EwxCmuKERX1L+RAoTjdNlNGs4PZg1l5CGdOWQ93cm
YD8v00qOQxQ87qivhRg+Fhm80Keo7jYokllJxlFfY5rj5EKB37PSGox9AozPRR+a82VD6enQjcSe
sb+zNCSAIA5AOqf/bQ/ru69fjnk2Z+GuWkVMDqrQw/dCYmq8Zo02c6LeEJDB5CYZWg1fKbA/WHnJ
ceLwrWmdd73bLMQWUh1hsnD057OPrzgGC/Owv2FUAim1ZqKAay4aa3RVqDmJ3fbexiWz/3ua61YS
7Q7Jx+xxr8qHqLh7wb0qdZv3py2wG9XzJvEVItY7uRLnRtPEHa7dKomv6YxcKOrRVjnrDI4adY34
1bNWfG5+fcTbV0gNyu28dMT/+B83sL2Q5Uq5NnV97WEOupr1qhba9tnbkPDBwxdbjekrRARQDyU0
ZZfyfUSwVX6vQpwKTONGNFZhhUQKH7wJwxs7UjJpUuhcftdcO0r+DJSTqIiL4DgEh4Zebkd/++hb
hW/922y79UN49daRwqtIKQGP1dXhbIpwecWlE7dwGpZUyNTbljuAVRSh/aJYWGFilorCsCH/XCoq
63i366bgJSqOQCJEwcrux0RCNWvs2VutgYvhDO0ebLcBkDWgEhqcIQ8uOu5ikaIELLJZ+Q1KdqzT
KgiuvKyMbyuybyTd3NoO5f8Zi0IH4B70sx+Nuvm1uazAjx2lkxhsn1uHhafga/RmFid0U+WiKa2Y
8fgPxI9rkFqKPdVmP/6xFobTwVTyKaj/qaJVJ9CD7OGgSsqby9crMy4mmhAgqvVbp6MAnUE8wyPH
VbNWv5jlVLViAFDRLtgBu9mIOZndJJnwqvjD8YiwFsm+p43J5ufsVoO1s8x8iZf5Q8XDnEyWVYiV
Jn/sF40HsC7vdi4CtL74rXG0f2x9Rr3UCjxfNLddLbf/PXMQTn+hu9+iv0e1TihxVITcdkfBU+ca
2pKaX65rHM8bP5x+MXphSDSeXmP0J7RrroXhFAqJqVRzqDJCqnFiBtH4c8GosKKaDsKj6P2nYWfS
RLJq9WE2hfaoyMwF6J0DGUuVOmi/Mb6j6t7fAp6TOaBUzasKXOR6BKk/ECssTdbGUax5BYG7m+/P
+WniuinqwfqPbOqQu5KstdVIA6a6LCFNNf0wt4xpQ29UeZ6q0+Z3Cjw5UpAb/tisMnaXyo8C9v9J
GAD48ehJkIfETvaK2lvj+fbXrHVNTB2Ikrq4ATwph8YjxGJJlyLsdnxjjwtO9nbtwcfo2nX4g6gg
iNVDUAV0GwQwycxdmxwvbOSLAvvyLxz/fcaWXp9uWFsRnjT6sBxpsmP/czPKg8/PBSjkoZBTmSsX
h2CcDb77t1L6NBw6rZKyCRFdv2Ze5QGxQLkn4URyveD2akVR/cc95qEtmDQ66lRcARDfdDTbuDy0
uRQ4tb3CHZwNt5m79odCJjLj0cLk9e0+5EeSZtiHOd9GCnrP3vaFzP1DNwghiqt7XaDRQeqY7SoS
ocXnz2A/8cFYB15B6d3pEDmQ/9rE2gQ+eW7RR2Tf//y1TXl6aYeDxFA/zwDEVAncO1IEIF06BnTS
ho9x53EY75BTIhZJ60oKsbzLGEE9WiGgEyc9IEk0DWgWbV0bODsUEUPQMF2MjkMV+rGHKKB1Rnee
hZLL+BLoqMDjBwS2WndVocj1FYdmn9H8bFDSaHrDM7tzyh/GC8neImWZ9Wlst0OjRYhvN3ZPFbGy
iSVYwQ0lzkNVSS8TKXu0heJa0d8MTtgU3JFKXlaY6HdLAM9d2KjT4i8Y9Q8JnZWqIGFAoGIRgwbB
ah3O7M/hL/zxJeyVkOJp2NoG5o93MXope+fcDZccIHbEux/JXidmPCxvfvV6NypS/sOVhppRtYEo
Zl8dq8ubsfFMz4qP3h24yNcLFc/fKxPXghS6YesNoyNDr0SRxbcQQ2i//s8EAO+TMzONIOYy+kLI
YKHcREGb07uHUTmlLV1z2vVCdwm8y+VNReTXGlg5j/65p0YoaHFMFv6XQ+hGdujqul9wUF6jaeyy
bARW+Y3a981WCjoxGHaE3RBdgjcZHMDeUOWchXQw7LkKUKM6kOdXQmP2Sm7oIDG3qs+SOwdCMVxa
mupnXDfi0xbR0YKBpApAt+qVfB9lHUXX8d88MrrF0DKKwUGwOVgErFNvSBY98YS24YZjpbtjR4yy
ts0ZPMP/SprvTO0eBqErQsgqpOr11QwN3AZWHLywYfDxmmlLHz4kpMVzanBbuoxcRabWE5JIsivQ
PSId2AV0jgQxu1JGPNdGPI0vUOK9J6quzl7JGzhwuAffUHJBrJwuAwiotg4THQJSAV3aK1VYEQbL
PXfbxCLMFd0Q1NAzxvryqXLNhtUEh4WI3gP3Diupf4hnLbZ5bBVEVLDGUAwrmBh3FTzLA+MLm4eU
uQJVGq5gZVjaRL/eIN97djd04tXJQGBO2ciBbrBeLA2InlR5wY7/F43Ln/en44EUY13yRln6Ig2l
xQjlcpuaPQZvCcMzHCeqe7HmGh2hIs7S2sSoUNiDdEM2vtlSFNo27F6BQx3I2n8oJfCgos41tr8x
DnwrPhxEQTAZjLEAlT8SQ0ZMHgk1fuVNgTxe5TsAtmmQQ7msS8/z5iE+MbBvITnlC1+uBC/3zMo3
4lMkzNBMgw+0J0EPbBdIAwIoPW3W5RqYu3FZCTpFZ1ck8PsX1eKhO1FVuaUOyZfWU1+ay7TzWtkF
vtdOw7FzGaKUaHCnz4+ip8cGI5ZQh0to3uE3Sbafg0IEjUoA5nZtHE3aIkc+j9S+qXtT7HT4uyPY
X9FvEGv36+AZppuql8nF98PSlCbZODGZlIHggnxTVAoItuiqbgOlWD+ZS0S4qjiUKILTmXNohKZw
MID10RQyLvCajvsqa/40izyFYs71job9/syPWmWEitJywg4hZ6gVzFOmqHfhvC7EbzNr/b+qHACE
sDqu/Q0UFRqBCuRinq8+E0xeI4sb7uAXQnrG8RlGd1GarDQcQkwaw9EXGj7f5DA7ZB3QqXLmVDDd
wZLjKjIRAmeBTAG5pIEJnToc+siw84rhuZmjtT5peUO81L7PxfvYqV+m5B0r/deQx2dZDCCmjnVu
ik24yhGF+Cic8Te0vu7W78K/8BeHzMxn3A2/EMuejK8yFsrvuyZSKQ7N5F6mEiNkDkHyMQLbXTn3
UiHU5Kl1Zb+xfbv50snImSAqRkDm9fLCFhvzBo4SFEmwaceyhnetoWm9KslSMsOXwKX5ar2ipefp
yHO5D3rBW7TvFkHEHiIy/e5Z7XezvX5uONWlagMNnr6bRUfvaeY/RW4hdHDmGZlg10g4X1hiQ3vz
dnggwPoKP9fXwClNawczkSYWc/WS8A1xQfpU4tAhkm9Fo80t3ofRM9cg+VT5jCsuTFAcsdqrS9tV
2qKUEtrXgiil9jY4F8IHwoKAtO6TiLl+42+LI5EKXdp2Z3JNmjUp+8fMeKJfUDFpi/JAxqyALYrx
+GUizW7MVwHwW6hu4SPk1KS67KRHIVhspRuSOxCQq9vl8bVQFUy6SWfrsnZ9mfI6BF76aT4ipie2
2gtZr9MeXet781gY0NKTKkxBDWsw1TxCS/Ila0bfka/rCkv5HrtvAgLp5PZCZ3vfu+onsfoivIyR
xnqP8XUD4zVqBNubkUAcAEE7ZdR8HQcx/e2HhhTOH6cHRwuPQ02cEtP08u7tCDZ1cIlctXoOLXEM
TPle3zRcrhV3OgEaE9o2U4Pil56pCYGEBHQ1t2NLzpBwAMxwjDC/8WkMGoIKFFkEqUif/UAdXLCp
QCObUrm9uwHSjsEClMKw7ot82cE9A8FuSmHQ+PfhGFnlbetKt2TVzpOCO7gmRACs0cszVPRzGnos
GUh24KaykHZ+q2t6K6LhdVe/cL8uhkGcQTQoN5IBKUwdc9Snoo9S1gLL9t6Fvd8qxlVibnMsiXk/
zxp4HPcUq4ZaLuLRqKJr0XcD6yj7ZPwLDxRCY1oSLbhaxyNwpLCpi22wCwOMRBT3dSxRhkQhkRan
r5dHbEkvLKk3/yNdQgf+e9frZUeUX7FSK0kcyA0fr1HpUdEehBtIUukvowowPktmJ996a/R3MBAW
ZK9f/0x78t9BM7xZ/p9qzbTTe9kVi/opQ1ZEDNbzoHDcAEbMLGmWRUmmtcAh9ZqKhj3mi6ncuL8y
NY1D5liiMgFxk59umxTc4PgSjC532HUR0x7R30IANHlhZ9ZDFgiF66Cb7PphkaRHB1Y59o7DUZrm
lAJ68kk0GrK/rcMo5/tD+sUKUUl61Vwgj3fib9Wtk550wUnzAOM5J9/NyU4gOZDQ/4A5IRwTctsW
RXNDpHkhfPGdMZneIV2PwSohjXRxwJRhYLDxKxLBCwHfD9WX/Nm7cZKhQuwVRQtthtf0dupamgQz
HV9vZ79maS68376fqMrsFGxB/pOg4ejz7XbTncvJ9UA0t3cYmUpBAEwYY4IuOCYjefBNDXvYmMeE
uoHKo1bE2SfY6Yen0SM59ap6+z87LO1+0o246fWnPcc5zs9IpbpFZaM7EbmiA2i9NgcpDGTLHOMf
zMyKa1wDPfGGi2Z594T7JJnGbMHwo2hsX0VHE/Ovql5oor2a+baln9h/gpxdMzS11605NXkc0BSS
kQ1kaktzfJAXleLTqwYJYSvLWRkFgzT5xT158iSFxUt0xK7NsQ1/uRatlrEs4T1ROpqv7LqQMSvx
3x+fbib2HeKCfbMNvv2uC6VLuO1nDZFN/O+m4wuwEvBwMCE9nR7adJihvjDc8sAEGTFPcIXL26O1
fsF4zyZJWoLqq5nc0rNc/mVopo9+61Mj70zZjU3tSS8MCQQ0s6CND24Fk+mKek14Dw2K8lfbcPBu
EWlGsMho7VbQAfWKxi/aOf/AuehdF1SIW2eIeIzUqBEZ+iszzKNBOF3f/RuVtk5hI/pQfhouINH5
JUtqRx+Zea2RambfwtH8uWo/EruVaN0toeVucuMWMuQPFaUaQm5Pql1Pw//t06BBFv2uCiKlTsXx
Ai2TUjJCpchnWGmuq+cFWbD9t4kqDyOLdkYhpItGkrwuy1AQaxTIZ7gUV9iyfdlwTy6Q+FPN0jiZ
xTD0qVH9iwkoyUA+PEz3Qvvn6G90b2q+Q7OgmCvBxqmdEV6/y8sZFYgQUAdQL2LicmaFiTuLTbLx
wSfdmzD/L4EhlgYqAuTSyVpQdl9gG37ejf5bI+dMGEvqBqvFborSQHJ19HgiQmUJ63fTBCrasESF
U7PQ2J98AkSjE2CFCY/ZvFFu/SPYg0mRRIpVSpcI46IpUZo9CIcqPS51dcyp8U2RVJs70lw5wW9N
iWHJ1XL+hoL8mEzrM7wfJXrukvMLn6DP3NTKhCTbIWCoWDOyyGYlT5OOGtYVlnxYbkP59/XHSgJt
ej5Xz/FxjVMau4DZEEr5KQk+xQynS8ILtraPc5sDP8HmbzqQC5SA2OOr+glRtHJFflprxbVwaQaK
V5DaS6WbSAelLBs7xhj7K2PDC+tUkU7gTNRBb0+eZ2g9UNxMPn1h+OIN5X/uPI5UmXH3ZDx3X7oU
9t4dqaItp1GEVAYfkKAOB5npeAM/Ap//K3prl53nn3CjzSDV1ppY/SfTeu2dv1kIsKa9pYLqYB8N
MVxyAyRW2b55PnZtG/EjgSe/bSmfm4LixyeLP7R7DPU/gmb4qxKDvfkQS03uxfkwrhz8aHtXimjX
d7n/eIvjhdcTmKcuaUCm7IeK5rM88oPkyNEfGBYPAH6y2eC7xFOqdfMn6d7+gfv9oO+1LlSrxFME
YLu3GGTczS9DoKpWsshw6dVmEWB/5g+gF3LiVadgYQFxUVgXcbTLhx2iYHlsHrCDnk10IB2aUYBk
e2vDOKOPFGEVaozV0OOo1+4uq0PjpNnKl+IKqIzJjmkiYvwPSaCVmrOhXe0LRkw1kCo9dmzH8b0j
g73jxe0/ojGJBfj79kYHMKS8MEULb9ho8JGOVORYVJdZZ7PCxritK0powxnhy++qL7A6G+zBpnYq
SikRuqQew2LfbjseYTYg3mwpXjoXUZpOKOZU0bEFC+iP50rEaLKFW7E58VmcSvPJqpzh2bwARE0d
eiQEiGCQgR6RZFcPitiS2XEaByZxThWBA2BCo6aXQj5jffes9Eqd0RwpN4y3cUvk+AcGfqzvSQR5
rbcOfMDiaox2Cz013MUV9jCtk0ccHY3htnMZHOI0snc8K0h3z01JlulSwAapqV2C6Ehr/m3BdZvn
0BXyCOsMwonZaYjlwy//HLrRVkzGt2GeLBlkfpOJCNAyRDJKU+Mbb6uUDNJ2OYTIk+Wya1FuedQt
cCTxm21zQHPqLdbwRC7qOqRxEAi4bBX2YLTZgZHUOe6OCHpGlvCqBXdAXXBsLq15ey01T5s8o+bk
d9zs0pASdzK+yPnhSH0kw1afYLyueRwk29hXp52MX8nCiz/3361CZKO6nKYYNziFsnHCEY3pbUmc
VzFCy7pMIrbvU0AloQjeQ+r86sFg8uBXc1xU7nEuN2hcFkABzQxG0VCu85fdFA/9kfIukv+AwHvA
6PF8P1a7fooduEgoLnueMY5dbttCGZZ+m9PZ9MQ8xAbJQxtxaRlveUXu6x61sd0KhYRVt+HGfvOQ
G1Ge7TxR9N5snM9zWP84+q5SwQjMECt3XlqvoqU1pwmvQ5Yz/8fX8TDxWe70GQmpvmIcS6A1bf/r
aV+BqFV2mhFQkyYAGZj9JhA5ZYYADvS9MQ2b0P36xbJ30Jz8TTk2da7N2qQvsZxrj+NrpPhujQpx
l4Z0rj3sPUahRABCmGgtCPZC1YnWMwPNbXaOYSmaorUxsmU0a1J58l+AawnZ9vKhGkLxXIXMcd1r
oQ9LYh+hPCg/+gaYHwOxExY32UTdawKMRbqsFioB+7ygtTuYzPG1I0UFzDl5FC23ZO+u3z9cUnSw
KzeA3CPMJd6UVNoaT87XB0wZ7dzEqB4QkROhyCWbKgjRo3yUnX87xZNh3I6UghH4m+TrAPBGlCWX
sCHBPFIFupTBh/51vZr9E8wnY2/SyJNOQDvBYOhzeVmA42UpOrVXJ172vDdzCSEAfkKFjRI+QtC6
8SPHQtwsipGFGWqxqnpW2Jl+VBUglnv2Qf77W87wQqLY8rp2ES5wRKuqUyH1eyje21iAv2AX+V7F
dFCwsk6XFOveeaAG64kRbhjszarSAA38PwxMGvZM/bEM/36WVq5Em/c+BibOcK6HyMSdRRZuMoYN
nIkVTS1neQH0hlsPBFvOPIkHOSzKF1JJNGIw2XFnalrDsXRx7TqK9r/3nwjmEOD9SbjQpPdzT5M8
5FbZlAzGibk705lM4VkfxOUi9o6/ZDVDimpPhCQmcUXF8SY5qtfQujhPdLeUV83fT/1eME4itbBH
cbOWhSJlc+ZDQvHgn/QHfEyw+Ylg0vpR2eTdrf7kmJZFW8N35/yRvALgaYAloC1KbiThrg1RQ4Pf
L/WmM9AQDkb3qdUNPUAbbhr2Q2sVrOy5XPKWPiH0RSrWv0+IWzFzl/3gwYKoTTm50z6Y8AdnU7Jv
KmtNTuq5JjjKJMh+ExParoTHnsIIj/beaSTa3cJp8NRqHvE/wRlsbDbrtNRyKafOLgiznuyhakme
+LQdos+Xb5e0aC5JTWMuvrjVEwIGpKJLFpAtea6jHhdmXg4B9CNCGm1bU1gfUnSdQ5nCmSWF64Po
30G638/O3RufYMliXDM1ApZY5ONouaZovIf//JeX9zXf/qDP5licRGGFrySK/eMsMdJLdvot2X8o
L9YUtmjtrVnm/LHggvwm7Avda/QDPFegYmYoxmAY8/WDts27TzRgw4oj4mV4TsUicr0eK6eNKF+S
IybKrG2RJ1YLLeK7McPw3v91cYV0xrmJ2Wypg5nXekoWVSGTioxpVRU/wZ+sqVQkGk6Gq0MLMkym
hQVTWgd1uGaY9CPqO9Y/WzKchcyS4AUi6qlBUIeZMmGFpcd5/6Tn13SIk/ZezKDj+y818Pss5nuC
Iy6ApVjdo7yePqEG4/p6t4w8WGQtWOfviOnxZ5Hxz0PmB+3z9cgewxTr2Un16Bt92sf7ZDy0n5db
OaWQNxK8tfKroPWTY3N01vWkSmgVZobibd2e6Fofb+9GcMorJtHWV6AMiyQoMFJTfY+G/2pA/bzK
h7MkJ+bZycOg5Om2c/3FHPxuq/HXHkW2gMnhPj3KNDBHV+57dg01mW4cSZiTaBbIAX5sY3inTCcv
Tz5g+BxGQ3eVj06Lxm+n6nV7RkopzqaA1G9Og7MC3gleCzQrjT2qOcgs4ffm/hewgWScRHctXluA
Ke4Er0X9QYdWVAZrKu8gUtVmmoEwHbeeO6nOqhnF+61a/jcKAuZ+R1xpV7eB721gnWQtRvGJ/IPC
XKznMdwZnz1zHH14Z5kyEfqQMG3qEG21NSifdL/hTZGJhigckwkjAele2LSJEviit5XoCUG2NSkU
cwVZqA+TXJly9/euVSaX296gbWu5hzDRO02YMN8E0jRg98OBtlMl2Fqh9P0QYGCwPHXSrNz4Fpu9
tfF46H9RW47kHm8BH//YNwhUnYBYTpng5BlpR98neLU3aBBdprp7H6tyFV5IN8/ryp5xDOFwQ0/3
kKfjiACRius5HW6O7q5mGsDQN9nkphvyXsSapBu7H0HWRLoPozTCjyofNsO+/Bq9ihPbaT3HpFBj
mUpYZTQ1Yo4mnf80C4kiRkP4CuEoUFJrRF21ztXlIVb2z0qyHbUjZsd/9B/5z0RefTH60M47FWET
97YQT0e5mJrsCh4dWd9ofMVLH7/bLn8QZiBXeA5dTlFKozC28V023JBEGXmUxHMF1XK8Yz3dg/I2
7L5vNMiXCFYruBQfUTDb04haKBoOd/2gdn5mnhDVgA16B4Q9OqRvHfSNnfNUQj9o4OiS4Zw8YCWI
nxrW1dLyjnXj1fDTiieuLYt32Epz8lpgZFVFeiFK/Lpnn4QqX0XuY+b1CX/6DdVNYvw8PHKYOcBo
nl0huatmjToViyxnRjfD25Ch/0iObWRAs7oTTOTsn8PGCwsKEExdFQNFOmEB21A+KvpJKXgmFct4
s4pmnvMRv8BMa7BgGnDI15kAk287loRelxBOSvNMuRPjq05lPcTBOymonMgoUx1FepX2sjkcq32C
gsWNs5v4BaNLwvMb9sqQERyLmiIBt1wV4sBohTiuQjwd0c6CCdSdC5AIiMparoqc7R1s7uYwiB1/
JvtiOmm6OtXpx8PXqZhyexefXYMgmps61vd55C2InyALhQMKL89r+ZKTqZ4iCSZrjqns+amY224S
zi4bS9DoRPP7qTRYNA0qyKYtMe+fyjQbxrfnqZyjlMh99BQks57mszpZ00xZ+JUbCYDm5yP6x8Pq
3GaGIdtdqMiHvks1CwfLQpDoTC/5+vlRM4jABd/0gS079Kb7o7aHNB2jl4YQN9E/0MWMUzx7GHBT
9i+4T388bhd8ZWgXTUoszIuNeBGPMvKPfaZEa4fsyQYBt9ylNdtcy8+2Fsuyp0VPrOzDY/G9/dhK
pnvvevJJuDpLtAin4Gd+wfGJiiRJSYCVda9BruEqaw6sAuSeTIWdyUk/UibRNy4Pa4vurx/oeXft
iuaVv5Pj+LnRvHeRQjrwd9/X4qdw0hN9R8yTqe+rELZz7P4k7u5XkaZoOtRpFIK8jPap0XGPdltL
W6WyepeA7X3rTSR9iDJmIHR+AaANbPT1aXFDJDhiB9cPP2XT/qFikOKBdAo3Dwu6o1oYSDRgSNS6
r5xsNK7LkG9+EBOisJ4fQ/LV6qSKdWj0TwnH1HXH8HfMNY3X0QyOefGg6ICo0YHwlcMdttsew4ca
RpNxRWPuTfKFLlN9T/Nxo0RRiWh5g+nWUDEaf7ksbqau2Nnu+gqtKWzD6QWM9pJW+5zCdg+skV90
aVuFoAEmez6tNEfvLkUVJNOE6MFuy5sFGv5nbHJddF1xEXioEb+bxtvnRyYf1FSe/Fdk4AQEV+Ok
8fhvz83VMpmuw15PRq7cPfvARHbhF7oaq5OBjhzHRlii7P8wpTIMyGZPDDJyC4ARnhQv/CdrGnN1
XYNGc2yGeKSRDCaHiPk6Aot+BP7MY1pcEzDzS4r1sOklv+6lDlsJv7kE1Ffuk7NmG/2VSs+ukYvg
j3mgOS3vgDjbU+4gukfz/AtHwm8Gpk+Tacpy3EKu/WWwo75aFjLmtFWOrrNyh0gItHtaFMf3YQ3Y
iQsj3Q03WVylxDDRWA5DhTcIxJuexb4UE/jzKLmdGvly3xNfpb/MPOnD4PiEG+7IWR3iXo/hZ4k1
u+l6b4ucUr106dDHkom1L1btq0g+QWn+DZKlCU6RixVHM+rvawfo9aofqR6hI5voRimUWXLTioE6
tjhHGhLXDNHwUB+m2rqc2+U8CUV6t2/Onjd/j7SRarthJnMuYEmomu2BSEYLl++N2CZWmd+feQ/T
BEnydeQ0B4vsmgMvGp/E1m2GiNgkJY0vngnZpVVkEzbfxnK9ydXFceLd+V8+DyzWJ7Uic7CWRI8h
H9NzoFJJsGigc6SQ/RMx/wQeyrYwr5jj0YySDvnALveeM+rrdL+DP4oRrW2e5OWikT09r42hsx3i
4fekhdfJgpzuqnvIPhAmGfqtah1z2t6sTeqa2ZELgP23jPlGFuG8kUSWCck9HigQFAKV5WKvCPzU
MWw7aI/3JuPQfnwXV4udWuv/DJVo7A8t9bOOwzTbtYKPP9ycCRbl3eqeNX0pQVOoeb1+W0v/coPK
kOUFykUk8nv/7e7tfDghS7TcmyTGsxhXoU1WZOcEhUjmcPzXJTTCnq0Mki+rp0RBQKDctCvrKbW8
54HlYz5Rdd1wIq+cF+wTZ+6oGHC5xAatk/saND3ofv6Mtuc4N8fGBPksz6QJWmJ4KxyG/M+6owi9
7YC+xTXah6oUMVR/kbbEx4jbmihhdBtqGGWPm7zods/GXBqDNP46MQvJxLTIctKlxw9colmrguFc
/aA+4rHHk9fjE6o9+JfiSo0DbQaJFGhunRss0r9nM1bnJ9RyQ+Yg3YuFN7qt4evWZHbuk8qZ/PL4
Tpk0yupaq1MPmoGL8jzCpqbY5kT5mkqaiIK1LGxJI+gwgipHnEDH7apsNDW8oHrNZXwwTBFnYaVb
Gv18viv4HYwapTaqe5qERd4XPZTV2cBMuLL1VsHqCjkMWD8to+8XFIjKDjYsYbUWkPklTRxel2k0
e/jTozo+3argTM2I53dmgl6GUnmPT7m/VNgiCcgCLK0xOTDyvev7+YNuxoNSq3Mv9TKreBY54jgB
lB9XO7932ykF9oxCI8LUrwZQ3JN/AMIdC60e2BpzapiZaTRm4d/dpBqB/BpXSZSxxs4KI0dMaNXc
Ix4eJpJRkugTKtzeKd3AP6XcqvHDQKu8tAmsDbCmNpUNVCInITQ7fscZxVQwL75jdq7jKQU/iQNY
kVDpG5wrP/aI+HhLBsFbhd2kNMlW+3ZxpTbupEEFQeJvZmLwrr5SwO1kWawnjbv8UJU9S3vN7UuC
eOeoqYnVH8TYNfPdoXLp+dGnj6PGQ863PLbuA45i5samPlCd/8rWf8FiM2zNBCd0eJYmqciuRxLT
hI03jTf12LWecEMcJkkETqqHqfkqulaJ1JnHNtm15qg5QHNMtcDre0NveVad+U7DIpABvJMBJFu2
m8cJM0kJKprWrUtxR1st4GtsMgTuHaC6fjJq42U/GMy3QZDvsi28S2aZztRJ9lZuFBTiA2/N0fV1
fC/OQL3KLxZzguwAH1pgM0mbPTp3afYEphK5PJwTfK92XKAHFV2bWwlsKz5r3hhF/Bh5t5mp8rNJ
qO+rWaQDQj0yE+1xVI9MJcXIxjdXsEyuIX1AFkZSTaWzeOduvviDKxyBSFOasg9pbw6h2jRKvNJN
XJhl6itJYmEMBbqT22WFLGdM646iFqkprD0QzzXVS4fImr/5C6WWnohpxutwWqdNmPdBt1JmI4JS
yZASwGwsJtjWgT0Xaxl5a3Q90lYyYTICB0TcsCXI4+6Pu643av6W7/n+Wd38Rg/bMw6ctXmesSfU
+21CNNyyeBuoEWSkgoCouLBUU9toJoUBHb9ebOZ07mbw4sU83ScEb5cr/z8XZDaFR27BCs5uqZTo
pz5VCCI7ssb84WJJ4JF8uCPm6HAwJZNXGowv1gbsWxFpdiBeSWaIKopS96mv7fQ+IdQscL/6ZOnO
/8EzF3qxvhyFbAKor6CQPC9IQxSqeEXsl2tshtkCBB7RvW/GYDneNkBEEFjUpay74PAhr6rxAbrC
s4am5uLAX6xvNmGpxCEqGqWghNEwcXpRYtC0TlJWGkQLpcwtI3C30hvZbaQQYtClF7opIPNC5Jxh
AdD3akcrJJUH4olcIOSknSGacIH0fj5aRgK/VkFQjD1XV1araUdsaCD+KQJ7zEJTIR6HjH1sbyu+
EaA2Wvae+38ebHjZV0FziSSmE3Q4p0Syz/FsgegUhGcaI/W6sQRDpyuCMAoK5UROa3qjwGfgjVGT
cXDGI/b9ST6QR1h/MdvmqQf35Ewhl7ZzxAqhNqsl2E9c7AuLAl8H/fSXCbr2s9weXA8ks7McxFfZ
qq9NNSS0qrN7rnaW6MUueE+WFX1gcSSurwIvVLXNaLl9GM53+wBEz8X6dlixjYvy5XvMTlns27i5
xulrgZsAhee/dJ1XfNgM46UBzUsCJWNnl8imcoU7ola6VysfrKKKAPuRopjUxWZuZLMxjjrAtpOM
2bA6W93LQDHRsCsYz5IovxfGiJqiIfVqd9bMvJsnirZt5uFEAxhPQV/UMh7Qkfq4CuoTuEFJW91Q
nCmq0rr0uQXRXMu5lkDYDw3kW7OW6VFCZ/NFkH0B4afF7xfDGkdMjMMdSAiHyG7A+nIuIgZKI0Mw
smKfhzN7VGaEKFHtHKurYpBCGcuO2B3jl5aeFnE7aWLj/n3zaVsqJDZcoZxRDzNbkp+A8JlOKegG
wXYaX7S4BGkPmNP0KhZgj7PvqunFspOOFZmPRpOMAx3St4zDQI79m3K2acfN2OeV+U1eBYOFY7xV
P3N3jZU69OOcLsVnHf9l3wDoxipBquIUNcJlhkqcwmz9cqo+5O3yKsWENb3Ho6VYH+BkBaEU/gKE
nGEFV15PjreH+F0IrAxDPcLcWJleUV4ieQJ3fjvq0+WeaV5IqJsU+jgGuG3A9+e/drI4mGyP5LE8
n9iLtIBnyS8X0jY9SOQxrJ42i7kCz+AmiDC/mdUBWnIVpyzl2GybgERBmoThlHdwdVDdQ8C65Qs6
7+PLMvisezPiVB7zk2sLSFbxAAsMn7S6tb/H+DMSwmqEV5xSmK9IC5ZEm8hn/hUnXEDOFa8uvq/H
X79LRShqaZ8aYDDJ+NS8fKOSfK+ho/1HkzExUR5Bd1P8WcaGH6nrceP7HPefY51RmV+ay9uZtcrq
Jf95uay3nVSS09HE8PZNGAa8QzN/EeXvlE0CqtxQ23kaJc6HSzufQ4Bl+3JCrXLwhZGxRCPfzstU
JOIafBFwRRKp3t/Ygrf+klOnBsrDtwSjSmWtEbUwJFQ7DhgkA5HgmKf6/WM2U1rrYTM7UMWgpFvu
Foog7lV+597vt64GuS1UI8eBvPLHz1MBn4gfYfhCCCkX7pEX6IcvPtpVXUdQSU6PI8Fq7t+kxUGI
2N66H0+FGmnPTbaCb9QQk58PZpy85r6Fp8uZl2pSOWN4ZoZOn6Ak2OwEcRQyOtcboW+YwWN8SrmY
BNXKE/nlkeQnAPIUBZuecL8YWp3ecvo1sAtz9i91bMpQ2LF/KxiWLFQT6onWNe7gnFyDKnH+h796
PKeEFQYgrv5GTfwQ4qM+RofItKtu4LrVILPE0afDP4oejX3STDndpSDawETm4NlbAzk+lb0Or5C1
i1pVvtRjQZGJ8/LrH3L9JDVQATj2Vc27qOgJgbWwBRElQgf7ddQZYmLBr/Ow3xSLREgyTfu6fPAb
FqRdEe/qU47PGH+wbIqu6OaFoUQ6gdEVHpd+/lOGCGFzl6W+tNte4+hk/15FL8URBMbh8ZZX5k+n
FnF89fsc5JiL3K5ioOEqL4llwtGzP5C5uLikslEezcH6XmkKHB+qz5EUjDLNw5/LdRCy1HDriPFM
6KVzOtBreowIDuBa04xWQLqE3VWlAFmgVRAB9e+ri0zgomNPodNItijj8PiqXcu+GWMX2qKWOhhK
dR/HXDioB3N1q2z/hCk6ToIP0Zc4NsvKNxuS4HAsf0knTn4PYQcEujYDZB5/ORIOAZnvgVcsdVA2
mrBayDz4eVzFS1AEQM/6DT5h9eHWOR1ZhCsSRgyrC9pOXXt1FMgj1X5ZkLkN55oyzkJILNpNqU3i
5DtbA4ruJ3H/gryNBnSkIKQrKAKImU2JzLkcme5z9q0K4ybiq5b5+BcwEPhr9MHHOZUNXZjWlY3f
7y/WUhzwvClVLrgDLEMboxoIDZf+QE6npf2OTWEDf1ix55eVSRpJ0VKZ8d262kKfVClRAN7JZZ3G
WZ5qu6P6QtThoF2YNn7kZBcs3MHSyMdp4luDgYhbMWkEwyJheBo6qffKOnRcCYbzAMwqrbrwzpI6
KADwFsEuxh6dhfiECb8w2DDYgzqMOcmXzreFNhvjVMGQ94pMMZJJS3HlZffkq1FSD9YD/8ZYVOgl
VOxqTRd/iYaNu+dsQaAcd4wCqXyVLP9qBi+Lxm85Mj4XkqjuOhdEr3SCDcKaNmF9q2W9O4/poU/n
Bbzr2SKJwa84zIkesBVN51nRUoixufpAzAAnROxwS7KnTjmBhD/Bwsactg5BOKolt8IpA6GyQdwQ
2cGGwEadhsnDBFQHwmlcb+A/geBcLfLVPMzuFr3GqNT+q82LxufE9/uK7IvO1ID+oMzucu+GHNLd
wfv2uuBdWJyXRciGJB0Nhl02d7J2o/BSq+K007sYUSuXgn4BWlpBFE25R9GNZpQBvub6+mlmp+GX
jqVspOg4i2Jsrz2ExldVmy6lXi53c2YHLX0Um6C6/1OlB4rZQFQ1G8zzv1P05ucWeM7bk6wBgbuI
47SEOkxRa2jo7lHOpu1kRvsPBMp60w0qycbWrz3gQsC62DySVyAhJPcYyYDIzxUxqj332qKBqf0o
2u3wJid+uAMYKqfT5wSv9l62d6+rtemFW4x1T9lNMa+g6tCFzir8sngaqgngB1VPFv6wrsvY6xzg
zDLum/W7HLu+EizvYVJlFlHSTIMjCU8QEulmiyidqMGLPZUQSWiEabXbZwugUlMYm4hL0paKO0w9
IWvcWOS6mEDeXws6+F33413vKYR3+cUErX8JO3mqVdqD9WjtXE3YqCyvGjtJ7gAc5kie+nCZjcAt
VNX/o9coWBIIXYt6MyBkxqT2NIbanijJdzIgfh7QZKn7oEdpb35zH0v4XeJdA/CYWwntmPOSZrC1
G7mNVphcNcDl2xfUj2IMt0PjuqJ0Pk1avLbtbJ4kP3XByemdL/rbppFZWXIO7OBMcJXU3m9fNPRP
xaeBkwdtkbU8rDsgl19eGyx1sRdAarPEr1Q5Tuax/NrD/mrQB3Ffjc3sMvraL3qtbwgbYV8Xt8DT
uFWiJJzlRYEM7D2sIVeH9rZ4lxde9FXgUpZMqz9RG0Bmiz/F15+Xxd+0jZdJgzqjFF62OSsM8Gvz
PkOD7tI8PsqjCdpkH3G7GKL3WmnsDGMMSbeeKiZ/ICNgldwXfBsap8ua4DATX02Q2/KmQFb+hiAq
pxDiNB/rg7SHuRemQ+9hNn/cyeLBywLk8sx3nczZxVYh5PHDCWIGgeMgZhwTGGzF43s+AZ/sI9vq
VFuNSYsJ245KVZj7JOcjF5EvMAOXWr3n6p7r/BUHSzhUmvW+Rl7rh1zVD2QSE/DVldWwwcrWpnzH
JghaxFL7XBJbZatWtZtmNw1G/TPcYGhP2uEmWpeMhKlz3RLiC+vErD1KktWgg+cmNa1qbF0rL5Xv
z6NysaRwTbwMO1PZ19ngQi6Pz311k+JE0Ylp7Z/FJlsE01XRPe/ndhp6aKnzi68Dw4DA39MGniah
h8ZyZFOloBOYrSxsqTqZfO3UjZSNqfVVXRF429bZcdsA7RA89xL8vlFU2k6ZK0BBiJg2NWXDDfkc
LlYtAtOWihoEnT0JXGqsx8tjucqjy+4Ykt6LuovSh9jgqNUBv04SL+t2tXDFR89k/bRIg/EKA2PT
mA5VS/LauRPWUsEguHGZJmAVewQMaMB4pkBGZfAHtJv/0uQKvcBNZ9zWnsYwVEFQ9tN6DaktTVjk
wck79++ux4GbMGEcl2ZTo5f91fQ/7u77SKq5aKEyMYgaUHOp4oKjiIO+gn7vCQLvlCk67RRToSOs
tmXePMTuOHBgo9hGSdlbF7muwqNprL5l49gASDgXZz6tDcVYIGltsTv8u73+DHLe8r6oSR91XT0D
w6RHdEt/d4xkjz7q6hzCq1wmhlaNmGzd4I09SyKaKLlA25mVTD4+crLa33ouRzBobNIy/8zn4OgA
+OVMSSOPK9onhegsByUTAoryqSRInyoBZXUmI0Vvu9f5OPxwLYBWdEcHbn9vTbYSt/BFlR9zW1Th
wsUD71LdjllctcLoFbZG322wkGyi8cNiStCGPcfPc1rkOVqEFBwo8aJWvz1Cx7lxsmXGYvyKSkIF
RxCSXL0bqnXm9xd82ixo7CmbrdTMTsD6Tfw6lxBAPMhgv+aKMQD/ncuaUJjQjEemouLOIlJ/kcZa
AqLDiWO14smgbkmtH5G2JoZu44tE0burtRq/cBL3Y0lp9f2bzUuyefX6jhsKupwcDTM+WjrmsThF
39jzD0TGSq7fRPbSDKo4b88iu7nSHZ9ISbUJY8BjcoEHfnnwHFKcwU8Z3MHB2pr8mnOneTA4Z9Wv
SQPqCiHh/a0suCBbNoL+xzVkathuJTTrK2n/wUswP3cn21YibuSN8cb7JY5ipiOOjoD7bPOLeCEI
UK5pwxXWF5HZtLArSfWrf47291SNvwzM3xJHBr7ACcSHrop/B47yrHUdFz5ghFhnfFP7hDgI/b6G
SIMEFH9ilqcmmwN2Tr41O+jddmp2U2fTrh3fBRbViag8KujDHDkcPjWzcfpDrpgBAUVOHgCgHDuR
R1pcqEnvWKIcJePwBSpOVP9KKAChjjZx2jXb6IhFrtX9h60O3Zp8APggcUFpRRCysoOvtYLWkYcu
hlgqYapRQNUN2rHGBe0uX3Q6+navbYMgfCjLWdOyGtCSE9uBiorYuWwgCPu1+EX1WK4/EQ1NTuZC
2XYz84VBtTYBzvYbubcP1io6z6aFIOSoHvDbkMysjz8rnLsnWQ5gB1xosAc7qAaCJW7pm9Efs+cI
ximU1OKeZLFEzOgIxQQlk63ud2TM9JVveqP6SnAdnYFksqrfy1sNfdOUlFUXEBJN7bMYQQVOrANj
EOYj/bTWHaK1frJ1jx4H40oM2xkbGt3ANrcVW7xiY3wltpbWybB+/2/u2Liz7kYRlG0WFLZ2HgtD
CjVI5qCPGTJNF2Jw3iTE1zoavLnQ9wDT+RHxfV/Nyvq9ABijPlCZpRmoK+CZRcb8VEniHiMRLtxi
K5aYFE0VdtSrodizzr8sj/DZBwvY6nQgUC4UAhWq6/u634cmcRfUodfftnMsMDB5dNYufTE3vkdP
DZza6t/ZQ8/xfnIAXhdiVWGWUQ9QXXhh/Y/EbFB3GvT6J/W+a3ubwiCSOuITyG1R3iGg1Vn4/M+U
SriBxoM0xLqSK4AElIQnTggNJy7eETOze/2oEszpNxZfUy9q2GYCRZSvuB93N5zG2J9NPJSxiUX7
p/cQuBN8JShdE3Ko9D4erhXe5QKRqNpNb7dQamR5EJqSxf3NIVsj7+WSDKF+q38Z7YcTb6AitF6u
zUuMvHgZg65vExZ+TJRtnd+JOM0F36Yn18x9H2Jad/p5WCzRdsoiTiKyMDD2bFAc8Aq9KuNtHBod
3ZiVHQ3JYouS1/JhlZ+C7fhaUmrWd14LrOQydTIT24Q1yQx8rhEakH5JMCTNw3IrF/oDYup/Jh3B
vn+5T0AAu9m8S2w+kq86FnjK99HQMXO4dZ/63mcRBXwBmWfIdQIy/7qGhFjyCoWBXFUyEIJv5fs9
pFQo+nkGeC4GK94K7JfhFQNmhp6qgajG+HwT9ZVBIZhoF3f4mYVsaPPH7nFloJsVP+f9GNHd22kf
HuOT58W+Bn3cVNsV1cxGY7ZMZailj9ouQHBs4arX5moejX9oJ1BcwFMFChOr8+Ezk8zCRCLIXxqO
9w98obOKsfnWlo684dEGhQehAoNoe5wjpbuy9mgAivp44PwOyBA7TzgwsFcqgQNRmt2AI2xuzliy
+lp9U/TIzsSaWUVC38g/TgSHctqOtA7+GinfAtGpZPXY3SxnQqQosLxWBLQO+WCAD3yJmjhripf0
M6vq9N99K1w+jadZGcWKNGuLCaTZ0H89yGImJ8eEaqlpDaNnQAOkuDz8mP42xBWdFtbjLvHCEjOv
ULCR7NH28XtP4Mlt7RAQZiSY9j0cEOjLPJG3lzBp9hnNfyDqLtlrhqd1J9WVJ+txA+/Cch5C2mS4
n355T+QHJbSksSiI1Q7zsCJU2KkmRBzG0YImZvvwd1OxR58ozCgHlQIBYP0FZ+LufULvysn0IXow
O6XendKKgxjPv0vhWsVUO2/ejVjmYJPKZ49PdGwoz2xeIPNUb4BcMUzTAAr/q9poG74M3c83KnDy
2nvcNNZ1HL9ywdhy7iyJmRH30qClMU/Fc9fS4UIe4F27jBqMlMsrwsR7ZAKJx9c14yyupJ6wWJ1R
qYM1gQc2H2VTOHMsHcDKuaXkYps48sfZB/GpvCId7rAyX5pHT2gZCElL0zUI060Y0Q8kMwUj9JAR
19mT3dj012UJUzbf9XTyDDNYj6OIK7yUm3ktKHnPVpKrCF2fiOWazn1maUwEdbgiPlnS/1357ZL9
Qifyinl9cdUR/XMOSEzsY3A7i/wls6fpDW0vUbTMKUYBUtxpM4iN8/PLmNzrgewPwMFGwFd51p5G
kjXHH+WnB3x/xRScu+FIpGSXjWn5ZznolnQTAWNtTPgIjIYtuHmZ4J3kenAbTAtdPlCM8ifLG4+5
zb62bcuC34axQTV7r+6Frs4g5Ol6za2Vmg6ARZGmOl8kYI/kg5TP4ZfEoqRh80opC720KSZjK8Yn
BsiqfFYGid8WnB6IAqPCEyG5xHr1myGqo+Om7542pmqRgboEwdIARCcgcFZPz7s18G9PGsrfI5qW
FUePpoB2d1C9hbblzsuHhjx0CAz6b10LJOt11BPr+Epf5oW8SGhlvJs3llTEFqidAbeBXZGApD5X
s7VOeN+JHjCxf7UuCkdmq+ybc985f5tJEIW3RTCwYj+XaC5ED12oMpl0xWZ9ht/njRnaH6ptw1KM
YPAOwh2OqGZdZlUjCx8yEz0en2ysmx2UldUdTgNJiIXOC1O8aUqQP+ney+ir+5cOhzO8Sekneb6O
nZkOv6R4BjB/7v/rmI/+QUQSn+UhaQF59ajBVZGPQImEgq7M8GGSDDzhoWcs05Dsozi0dWx1LLuh
n955mc6RmKJe0dJPoZF+499/L0jrWvnuHiPlfXcXKV9c6p658XLllgPlELMHA7IWTLUbK7vE/N3h
TARox+7VykEVet88oFbn/PbIkP76ZI8TWi/DHPFBk1NqgymUfgQlXERQ/T3h0kWKdOfCogmDjM17
eFbp54x+TN0gnF9NPpacwxtcdDZoO1JkfEmO3q2FAdH9af8YGbplsmAkcyknuoekXnytfaitQUmq
WAU3Ur9Kb1uyCQA7dLY9/soqU6eJFVDLH+1hh54LByfNnKLuZacjsUkKu4CvjhsTq/15Wk6klnfn
3Q5oBukhSRIgy6+SPEdBkffV021vj4Y9rnTNQzDD01GAd/zI6dm35VtSn8ZVmsU2Z3CT3kbsdo6n
a9yPdlp8H7pJeEh4jlr836Kj2McxPlmi5SCrwqxIf030DyAxzx4jWOg2bZxArdT5D+i6V6hAuiCz
DDsvObuT7mk43wkWUfXmVqfH1sovH4+BWMDTcj6Z4pkQE0ECcyk6ICNdkUVm2zC6/HZtVVoNEVNH
YisE2m+4Upz5np2Z1NeZ5BxzMxpylN8ai1OhfpLpk59X1MuxGYXUPe29VfQSSIOvjCfeyt5MVim4
y0xqlI342q9Yh1MHlphnyWMDQZh3rr6FNOANhiUE57izq6bWbQUv8DDub5MCqeQEJYf7KMFz1VgT
Xh1xaWUFmhKhY1s6x4XJJZAhwgKReIwlk2A+lOpO15S0UaW5CDZlKeg7AMwefCgRpNAyYcrAntju
0VUcb1224cTuis2LgMTVudvfFQRmsClWouXlXjXTGwxy24J56E8uaVma4qH7VXlKPrpqTDo2yWeb
uNidEn0UomGZa0gSiVYlHu7Ttjmdlq0rkL26gNYajwOCbEpJDcQjoIehpd86HLHe+sw2gghIaLB1
SHmYn/8QEfwQhSPTfM/ZbLf8OSIe89oQvVGqX6ZvuBpmnJ33ahqIY1oTVIl2BDli74I5xEkblMSN
y52233TvwnbCaQ8qTCMpq0Qe55JK0TRtcVxKgEL0liucHYFRrAOTcOQ68LyzkNZ40ncSKiqBFR6P
WwDtfiQdrNv2yTiu/ufBU96s/VpriI0AsUgERhGP5L6KSPEtjmh8CTUWbdPJfEnn384vC4ScDJZI
pHXcU4C/1BtgzBMZ3xx+hGv2H8XWu/8jgZtSs0QWvK+rKFAxgp9lR0CyyDekJWMuFU78GTUoNZtB
tF+F2MGe9+XsiukrwZXvxtIPdVgW588eOs8Hpv+KGx8/31A8Km/k3OzlR8FOf+Wm4/3iLC9SWAUY
SLmJWzM8SJeHfugIfkiovxMU4AV+oeSoidvQDsJ+0PalgfiANe4SvR/kLuJbVcPEy1gXTkvPG93o
cA50PPMlqL0Hn1dcvpN79HyWTMS36+ETZXWEEoXlnIGJ7PCDvz4F7BTM1IFxekXpWZ6tMx1+NmiJ
oyY66LqCyNVSJScAmrZiUOcuYCccB4UlfbPLmjAPTTk4PPoQal2Od1fLw0aadO1DOw8LK8XD03Up
bY2CfRlwMFl2IslIjhiqBwOW0Cdfi+jQ702oJ31UXrCSASpYWTtdTT36Z7QrzHzb7K6s0TDPN/8J
HGaoXbqjEtYXsPZ6etkZzNZ+X7WXpC1HSm8MyXTKK56n62byZUBaUD1n6nbiaBhWVZeXNf4EfL5z
7cJJN0q720rdvDizHWCo8Lu2n7ZlhlenREnjQ0q6vfokblp3sxiRhkEuUhJYfawj5SVB6eC6o+r2
k91t6+ZIlbg5M9r/48RRmcsFAIK+vq1W6oWwutuZEeePXYxh3G9e45LdTPvpmrytInULa7fqvnIJ
cLl+/eMed38tkaR9pO472eScqO4iV1yNBEAdyDKSh8PuspF71gLd//zVWM8DjDinO7ItZfowqIXP
lGLo1sy9wBjZQE7oj4kedvWzIRYU7fjaVgixS457p2Zam+oU57PKbnTqAna2+jQ0sjzDNN5B78xH
Ow/oCm3DIbsd7i0tnv8McxPXzHiT2qBWJcDyFhz54G5ZYASzXSOpFiFTCnZlmhWf/vmhvTy1C+wC
oVdxQ6IEApR630crsRlsmV40383Qz4qk3W+kJ9f8t0N4t65I3G2LntGr8XYROkcW+Nh/owNLPGIN
Rg4QvcE6NBkVPyMvCdHvXVjQsjnNo81cjfBA1HpaSdXI1Q0JMy0A0EeDtK3178tO5kaoNNSTVi4J
YyV6uP1HRquH99sM4DxR1kWgEYB35FYLJJm7ypyGpfDp/zzVSQiQTMWsW/ENZ9RgheyeWeiH6MWt
I4ZjhMBuu7TJmKKeBAzbUpuWuT/B7gSGTaBIqKIKfPsbJzULArdoL98Nlb0xSFEei4CHdnGuSDiX
OSeZY2a+ifHRr26I72wvRt8SBrL8OxbR+dH0+sa0KdeSwnaDTs+6poMx1susqtZ/KttIX6UwB7fm
xYndZ0qzWCVtxD14whchmNS3AFFL5ht/LA+vy5EZZmTDH34OZRKYB5qtO7SAypH+uqusY9Rxzw3E
hYL3wjdediFM04wggo/ZLFx3bYXQS15mXb0JZird7fYiAwAckbLkH3S8/r1XsSC7Y5NYGWPJ8wXM
u/yEz4On6DQiUw+Or3AIr9Nvih14X046jJFAYY5qofmUFpLpS69tgRQi4Tklcz4fEjikVWcrmqDR
IVUIOUpLV7Meeck8SPK4OKfjEgfpfiV/iMB56giWpNO/byFPJQinSuHI5xKyvHM+8AxGrgLJR6r8
ic3YYCDXos/TmYCfVsVpeXVbdtAC0zTJZaHT0KZvC/AOR8SKDxh4MwJEWaEOSb+3UapR/EKYAn/X
DXErac0I7xBlv55HckdsW5Jm97z3sJvJ3nn+tZIsGPb6UJV5iPQDiMHpdAeOBFSpDlfcH3k5H48w
RPsK11KsJb3dG6jBZPbzAFmSBRFGjnYS51jp0Nafl0Q1AWgds28gte6gPD3ywc1h0SsAXfJDZjCM
2nCxrcsLs5QtWKSDel035yJV4OeO6IKVp8B0lMtWk6iBBxjPq75i1sQsUHEt+shLFlsJ/7QCicK9
ORxBCnuKKmfqoGuEK4raxLFT2y/Sk+2ROdLxnNlenoVXtmjkDN2WgX8UBuexKiRdU1a9oUTWUPRM
DHKUhj2RQFruqKa1lqMzfwJpYr/HjRkRXCkC40e3puYByCKE3KNsrpQG4LrNwKSDLHs8QHFsiBbt
w43bl8A6bU47DHilVAwWZl3sMLMOK1FFjf5NbKWGVo621JFdvz8IQuBh+FBHmOm2+6W3rMTYUDyF
mKRTz56dT9C1tRewI9DR10mvfIwzIaPVxdkVLWlkiln6LjFi3c+tvdYSzaDE3+5dkmXrENB5yqgF
XVSqlxZH7ftuQ1YkiquW5NX1Cn/oLR14Tiz7850es/b9Vt6BeLHa6S0OvLiltwvcIL/cxN0xOdHF
xFx+M9xEK/imK0p/vOn7eVzwkc421exbXWulXW0YDdBf45Ucf4FeGgEX2klR8jnN+2RXOJf9bfOd
Lsl92sWgCGItOdOtH9nEPYC/AjS1NSzbQb4GtRKtZLBhL6vZSBjxxXwBlphk3YApI9eDh/zL2NAd
afdo4KTu/yCA5O49lLxaqm5fKDGreyeoqrtQmM0fPlNx/KWyUgaYyYklE+jdzJrqT3vpUN57DnC7
gY9SjWQyjeivu7r2QpgQc9dWOMFR+XrUofkkS9FDsT6z/Btyoe7mNk2BtA+sPKOZzfvbj3qH5Ojm
51ND0oaBcb+zCexpiPcYUzEnyOnbWicz3btyTpNtDO1PFWNiR5bjORToIWWvqngYe8RZgM8lDPYI
zCpHUTha0omfajR0XZTMGD9d4aydaM76JiOv4Tc5CoywoFuuiQ2CoODUQmn5eVekDheTpITxxbvw
iIUJWv2fxwWhS/z0ZrfUs3cwFVz6eD2zQU2UXlIYdnEOxiuVOZz6/7mOGzxYg1oX0WMZphpgbeMR
JneXX72t8kssHTltnMkgU16AGajyj2/RvyF/UJ0FWIJcShV+XmKsoJkasxcRtoKZtRg7ikAK5RNU
huWFfCMg/yAGcnK0eOj5+axKz6dn0paYOW3GvQuFoEX9WVKBEXhQTYMyhov5aMBpTSO5LS5qvrfN
ITaICuSAExYn25K8qbLQ4nbiF7wuHCylePC8C6u+y5IIDmy75BAOcs+0+1EOx8Ye88jCgMSztvdx
Jbbh5cdae+nhw2GBoQVMgHy96woyXA0R4pi4Vls2nV93MnlUXDQ1hFdAF4HOVGzastyYmPr+q7zA
1FSCk1oF9OWSlMqEppmGa95DWh9PlQ5+GvnRaBsVlFAD6n//x1ToR4cF7hPOz1ehKB+3q5RtzVs2
REpDBjUiE4NRbkK91lqc8paIp7A1dH18hBLK5LLB4JhghOKuDdB1E8oB8QBsXUXFEA9Xxz/+92JR
00t1leid3pHwSyhNf4jajqPV5RuV4gr1qCXkUJ8Y+juf73T5gyMTrdK3JG1on5+Q465a17QogaUf
WWAP0J56Nf2Va3ZbqOAV+nuJcM4L+dYFvqMba5UkRJQgW4uI0JfBdXG93yMElrOewySgRYVbGtkr
U0Lh9J8WGKknJgBcCXVI6/pVTSQl8jCrengic9okEnbK5zXP0N6rCLEZE3q26kAM9oPX2sc8DRZz
3QYf0g71KKT+j3G+kMIeBjo02ne9ewpOc21bqqp4k3AIK2bMFQeT3UZSFFPoP2T49amKzMmEIIQ2
STCtogulKkt1Kn1nPgrmbNQJx9ktoHxlakukC0gJojWQ736BOHin1ocpBpa0IiAYPFG9uiXbby+m
FMochbHHPfmF6X3a8BXRYs0/IQcea6SbFNpLTlYifS7vyXngRjHkPpfzVX2KXWOEC3hrvbnsDj5Q
uiiR2rcmyxvWpMlzsGuKjSEDlPH+qwKR1H7Vtz0PIgCFyDrWbiUIW77VaVfK8W6cwYyM+uO1vHjB
knMMHqXlUXwIb1/kejLxv1WaNTdu1EtIywIZ7qPe6giDrlX77EAM+mcvRTSAN5fVrpr5gzxPQ31m
KLs3Q0BlPxfMv5nv0ZDLP5+iuVSsZacabStTxOzSFSXiKul+h/YFKtibayFraVx9FxXYLibs4xM9
mw0r4AeZXFdD+97ZD8+3emdz7p8eYy/yZ/GvpIeTIsSzq/aDR72h2QnChRveaDqnR2QJxGY3coOd
ecU56c4ijHgSvL8N7hG7qFi/OyJ1PyOtD1xiB8UyFF4FmTvFP13+NnZ2GjxuBbaqx4FriWMK69kB
nqfzkw+C401TiMJPqYaODrBP1DAOmSJGpR05nijp6DLaax7fVjItsDUABp2FAr9E6+dptDfSSSPm
HTS2cWSaT/CdRIom4m/FTy3WkFeWuFwWSUbh9RozsNEwCbUd9um7qVe/yahXdNaj0UezERQQyX9H
huDFUUqBv/N62JK6OF+hT9D4Q3ISdki13LwYxs1lXRhnexqsZlW+JYgl/1YUSPqkURvLhkUAWwkx
l6LKpnMZ+asIYIshKEkb9i/gpXpxorPGeQC0re4XKZhMpvNRcoVF+pW4pssYHh4XqHYtUoOGj6p8
tFepNR1Y7e5cqgr5zgVD9vBadHAVvOdoAhX4JHo42lbmE8wDpT1HVb1dryO+vPr/dWy5pVPOiDSg
h3ceLLId+M592D1e471Z4Crd2VQeCmx7/IYmcv5bxqxJbwb68T9LC8XcVWP8BoV8TO1SuT9lAMRa
8GTSYuy+Mbpu63C4NTnY7JugBM2vPehcJqDVNVGa/yKJFO5rzOq2Cr4HyepecbA+99jK8ElvAnH+
9VwxU7KRlgoNqZHbaBOUIcOjAEifbVcIeI2GTpGqlix6gmtzNjFl12Nu18sot664M4tQAK44kml2
elk+8JRCTffEzptzE1MDO3+OJL1SVb9SK2hToB86r43U+VhQEys257dZ3d+yxEoYl8hW0jn7lFQy
YGv15Z7w2kNV1M7O7fTS28uPsLkxis5M6LUSEcxDm3Ho8DPgYG79nGzi8xCgpA9ERxtNP4uo+y+6
W+JmqWN1V1wiRtSG6+mGJFqOIipbv8mzHBq9ZJEboSuPnBJ+RRK/pRoTFiS2l1IHa2i9HORaMeCl
5/+nZ3T6ut6Kx7TYuIRIJlDgZQFTjpLfXZXVd6F8ctp+1Hl8cwDg+/QlzeAqjylFN6KXVaO65m/y
BrxbhrPDwHZDOJG0GolzyqGWmN8jIqpbfnf0Z3wSkp61uCWzdrvSqZGLjUWvoJh+uS2z4Vgbo44F
ePc4Viy5bQ8+l+C06beZtTSxCZRn3BCI3cl0jXyX9qzGDenXdeQMEp7PrORRUda+iKEYMacfShQx
b3gkGw2suM9whcndVmvrQTOocwoiJmRXgfh0L07oF5sjR9vAMmvIFlVxOPri5bH4JtbnJm5E3OhZ
xkMSzqO6g9xaeaUwmAq7M1rfXsSzYNmp9H78cZD3vIOczMG+0lFDrY6mM2wr8gxUm5Go1wsQDoZR
qabMMcb1vfaQblbg1yDXX+ptdS6kYzJJ/J4WJNgkuuJ3JANmAkHSKCtvtEzwSBRU/A+o/veqWAn1
Q8RTHID6gaifxRuNKJVOUW36kM3+602sAtTrV8SBavpLjL7R2gw9KbR7vWFKV1bWHhPqH5ihLyWI
a73vfDddy192amVCJ2Hd1dlu0gHjONu+giP5dAwi5eY6KCtGN31+BCaQYy5yfD4knCXZpwV8t5Cw
VUnPVOI8dJ5rhs1v6gWB459zuY1UUDZSXzrTEaMfg5y8PXXvZebOuOLyhmsRh74cERy7bzRjdtO0
m4VKhk1LHpKxXmI3H3zn2rbVb54h1cIQOfdgTnKLeOjsX84o6cMkZYZbKQEnpBVE00pnRz3guLJ4
vpNgYdwZNMcGx3f/+rFdgN/PM6hfgJajPxBeNK5Y0rolpYe5atc8mI5WrAUq1isffJ5GljyCXD1N
FRdzzVZmMmp2wfXdfC2mqKMUzhMbXksdYoKF7N7foLBxgy2i3LHc5SdPyAUHjfB/gteFqiXAuOyN
zEZDBgE0/yOB9lsG40Ox3AwlwpHZJog/lmdhIkp68LZ7Ox6jQ0YgQamJffq2bQNlu+i09LglGXlD
QBVzs7nsrTfO7kWTxeVz/VgLd0Xrpe6scY8r+9KPiMmNlOedFWlc9X/C7JzJwtz+WmYfdcNIdcUb
G1Vkn/1fkm/3v1rtqjO0r76OIpjOgOJfunkvp8w2Hn4SV2e7T8lao2AYqc5zP7ZC5UN/CYNjB0o1
B8M0d2pJ/nb11F4gvwMHUnv/HA8wYgDlrC20tbn76l+fyZcFiXI54NMujvBdY2UQTLYxxusp2Ur0
mfTEHMhTnLhVaKX12VBGS4kD1n7t0AVsncu7vMa9Ah+EGLi5Qba0lsqX3JWQI8bXeoJyMoAsgz1B
vvBxZuKrjR4prG8wiBV6KkRlegmrZh44YazYmoLtIuwMi1z2q20YcRcfuG+ja/3pHAzZzUMs6G3P
Ce4AKtNCY6bn4oXOhlQfkVzIYw9iLOrmRaA8GSNDPZLKijgfMXElXH3WEmkDgIEKsVji0ENb/7RN
glAfJah5oIPD3hIZwUycxocjpMwPKg0em2i/hrtSWQKBGcBu43Fl4sfvgfge/hSG4oH1rq41O/wx
/jWTJFIfZZz3YupTbkdT8BJXsyBB5OCmLqV6iDS9LpGnC3+TGK0EQDx0+vNErkzzUxYP3zZnt5fQ
u12hbFNQIc3No6R65vuHjksotskEMUEtUcQi4JuFWEJjNxbSmo2h2GnuSMNTIcVPrWZX5CST3f6F
GvoDmlqs+pzQ4DSVOImxGpJqx1skQnZhOMJtk6i6k32iGyxN6O0IRL4M/G3rkeUuLHivP1/ZsNkG
oj1geJmX43hy1EAy8yqlFL7tfHP3uD62yTVzf17bSmBw7zPbWh3HkIGVJsAZsyjCx2snWt1AQ1aP
aVbdJi+n2qqJTEGveroCbUKvhUWxZFaKf5C5AtLbgMGtph2548krzEcVUl+r1IMtJtHouGuPkyWF
FWUEMMPnBjWoIC8ifzHYALgmVr4BRhuN/vMa2UhAfOUTaZNopFxoDmeYZR6vqdf94cFy7VACOAUh
EB6WVikXdUyBKnVL1RfuuA5nrAxW/8O/2X5sFiQsRVP+IV3DH0UTu+mimcfccR872bFpPEhKtRcY
kQLH9/xo3atBjS4S99LUGFdSHsjB0cB6EavJszU0GmHwe6rzvuq9XAhgycXrrVuYWhA/EY8S0qBu
vQIRmGgvZtP4h6cXtkqlnB5NzkPvFZyMB4BbGjOskg6s8XhIZDSk+PyqN85eo9OJTxIFIiwjyov5
RxEO3BUTLA4ynjcdrtGaFJg4oOj/eFwuqZmxfUjZR89ZZtCSwrS6cgwLJA1Atx6sTXfI95m24+tn
cdtqFGMfyP0lANrGUMTdt8A4m5/3erLrTXZGzSdSfKgHpG4Vo6W3bPr266h8ZGust4XGktlqVKIh
uD65FCzfzy0a+TCfjrM738zWv7CLA4f8j6kT7mmhXJlQAEZqFCZiBVZXT3eCUynpyxDnTPWcXFZx
LawcBN5/M+/1LFUz+fVcSIZpLny7GvUSyOVS72TWuRzBSw4Rp2mSbuqKKLuK7Z57P8uhlHckhR5S
wXI4133TVsWfy3j0kdNSzAQWyJ+mR63d289KkUCjpGIcq5TR8q5p7ZKaoxWfPB2KUUHXefbESryi
vKu4HyoiQ7wm5nsKC5azNdtMPaQKw4g5DWlKBxREX3XDfjxKp9ZIugfpuF1HlXbn7DU4UwhC9XUq
1PbQYb2QwkoWjfImjRpVlYLW5gBEaEdHpwpNhfdLHgAC/gkq0kR+Npe7xS5jdOgzhVnXCjNciVtB
+U0poblBvvTvXv3ytmvlNo7pP/2tGNhuO5SdndsJBF+dWiZ2ZUtiJSUoI8e/Or1MigmwR1/9ktIy
UNQQN7i3fURCukKvXTyHQELAkLeFE3yElI+INYALYCvjNx2+kOKQDdcVFyFZb8q2G+oNAJbDH3ns
D/cbk+c3QJ1g0mbp1meFhL30sGETg2EO18CF2lh5xtt05VfEipTWgxeRQ6Pjz+Am+NsX1U7g3Fhy
GXPIMshZxUPs+8UaguAgsifw3HHClUltMGM8mAFf9ZlXEZwdvStqODtXdnHJhdkG85WQuU0xh5LE
bHXqYGJVrkhHWs2klZ8DydnBqnb4vfrQ7LO0saw+q4/MHqAaoUjKh84vue+Aw9XiqBWhY6fMTxx5
5vYL5APZQmY8M0Rsf0u7S7Q/lhQQjoyuIPNdIreX0+L6m9EH63g9+AK3ZvmxYgAmdb49G1DsMDDl
pD+edzdLaYoWRFRHgetSZn14Y9XlVAAJeqppJ9liz31prdZlMzBuRvx2UIyX5AZUdVkDPxqoTUTB
tG3CQlCAw5MA1VoXMuYMDFcGWQws9CLQC0UW1c2DThfzh2DEigV8zc9BTbIWr1le/S+vO5ccSnQt
0k+voB049xfXrfBf8Y0pFb7F1mDPunvxjLzqWTqibGh0COCU2bSb53LJdU+saW2m3jfDhmulAOJ2
2b16XavkbhG/djGYb/0OVCHlynDRgEEFmHT9Xd0Anuj87tmiyhJTSWN/dt647e2JBFH08l4oHPTa
NGeGWhFJEMx8RULIdItA+KRNEY9MfbvietwYLj7seWrKuQBBi1wWx/LlbVYGpw40FIqW9y3ZMajW
yXGLIaXuT43sPIkZiiHKmhJrQlM/oKigFKBP2528O2J0PthVkbFjGBYlqn2Ug7ixqMa7mVkeBGdG
a6ZANRtPfjghM4jJyqd88pB69uKxKBpr9v9kmntIwCEhPcLIAMalJjKI//n676/x5iudDloHATK3
P8Ylt3WwaixcAf0tLVQfeExvKpavK7aEVXjZbboPO+mdDOAoGaIBPQmSGkjtriD0RU0keTNX2fRW
Ou4/2d+Vb2VsQPEUBAIOYhUFj7MypZyP1d9K6uOZjPk2gHuW60XuSaWwE62S28gmm4YbrLdGyLs8
gnEIKk+eKeuYxup4Bfd9bqwMtbtX4HWrt/poxU4y4J/KIjevyQ+09PSiSRdDYy0PZ2puIRNxuEzJ
JvPSeZtz4yxSTj7B0oIwNeZRFUJWvBGGIr0CdC21NuTqEENk4k6gXF3aPAGeudOCO/3WzBUZuyn6
SiFx1fwlvugRdkb/ijS8d011TCczR7u9UH/T09VnfNCPP3cKJGFKsoXXtfnxlYpLQW/bjldA0XBX
QM8mW45QLtUmtyIyRAucy7ByE6l6DXg7+4kQ+iii82Qub0fv7kWG+kKMY/0WdPcI4JDZgVhrda2y
okJPBuGCc57F0+1WUMTATtQGOE6DN3LVBsUfXY52Kylm1Ch9cew8/oMD8hVTMIN6G4qiCKGIWcss
Z0Oo2gOJFA+JTJCw5Rphflun/ODp61bNPXd5wxFNseXtJNuIKbb5NSlbpho+4UOBRVIBlBPrnc19
uYXvlGxpxb1OLu9g7LTjD6wnv3H0ze+hQenpUujfhw6i8msJMa3kBWjdyA9qxxeeOZZDCFyl5Tv+
Hcvwyaaqf33GWTjHwEHQoI/B/eRCB2q6x+lcMw8+/+QCgbH06OEnFGnwwjg+zNMPDP4XpeD8Hw+X
Wt0Veh8a2Lj6J2xZrq+7rUZmWNFmLhxQ923hzO2rsDMYexfZsW9+GqhuQ+e1o2BpYDuE/ero9w6t
mLR+ea5eTHOGMw29JA4BMHVvIJLWjZjS6MNUC3mi8pJNS+2JK4qkn0OHtOGvsIzmcLoT5GxO7gfy
6dfu4P+9BzhNTdY5EjGSGSIFSrreZ4su0KyT5Bwc9KYBzPe7//aUm2eKUU68NIlUWOPlvxp4jek8
I2E+Q2a43MBJAGL2QyIxGpvR8W0EeQyWo5B84iKGUHv+yzoYOEg+W81rkPcEz7xk7pVEVY1gcp9o
HUeIV7QD8ZfPNVqtFm6Gl6w84XKMKsAgGC3j60zUTmypLwOYuNTi0J2wQkhSJZqXTpXgEmmZ9ys2
Bu2iygRXaI1f2WXa7fk1AltY1x7FLE9anuhCLnNCL+Q9qaqphk1CIbBDwxQOGyBrJOiRY8N6omea
3c429R5O8XHTYSv6QSmmRLAzKILVwAeNaKaLwtC4lX9uT3AXJ5V0It15C2w7ogbM98wPiAznYj4x
dy9R7OET2g9DZ8g8zrqPmJ6E1QIcHXDGsSth67CQZWyUGA+eeDOvf6wSx/dgLgf+16cyXgOaa2fp
V5jA4HX3oL6EyDwwkXWJ1fcZe2JIRMpHfSaPB6BlMDqhlyNZ8/tGVBoq+JF6EnaVav1wFHnQDpRA
XCF6eHttsWFFhhAdnwHZHwQn1KYhm4qy3jQXPnyirUYXnIUJojUlGQTGP40CaSkkuX0Al7E8EkQl
Y+O9wUimfPIq8sjjuKv3LYO3XSzigtzxE4ZaDk61Axh3qSY2OUNouz6DXQdj+IJgxDlkCq1qRSwh
tSRF5Y5y3sGAg92rCRSFVRgozxLRCrYmVUpBMDm8zG0YXrANzFGcHbIn5auxNvoehZ1pIch/K3jm
wunpmA481D8A0bH33Cdll/Oy6bTuLcH9iu266jDCh9+MmrTfpzIRoiLuxKPW4r7tfwb2pkAa8DtC
vmTU/KSDNCK1c8VOPCDPbvCfeTJZS6SWrJ2i6PD69KhTtfSWahumZFF8aaIESsazM/QyBcu4glWo
Hx77WPi4vB0fylILJMdnnBfyXbXpTG4l5DF6hTH2H/rLWFjsDOO9PVL6rLak7XxKHzKvlIKwh4CQ
tVcyJ2s2wUie0uZZ0ZJEXcAcJc1psnQXG+NfdNtTwHlLulcrWPKGPaH9dZbRCXlWmSpQvLHM/1cq
/qv1ySsk+sQtZQjEYzdBtOoWyLNz10G0TqHUAhzXqZspWMbTm0Z7ho5aj4H5oVdnEcZ86YsiOd6U
MUTfjpJU0xOayMGLi4tNLVgmxnbBiVNN2QWweXBuHQRH5KAGKrmBuZBLdjfrq06pgBlPkJVwdaAH
EbIDodpnuEoWZSIJWqwNhGql6PTlXhjfgRTEsL3kkYfanxZzxTQDDYU6Ao5+Un9AcZpn8AQrOsJS
9hhGL33ynJx/zLoUxSQMdPGrm9fO4hW2wv7m3t7JRmlWBMBFN0aNC3P5spp8UnGKZXWvVS62B1Kt
idlShTJT23j6BORRoamg8yjl6GHRrbBuCtCr5vmVXEVxyNbm9smgBlWaGeCROm79hRCz9kJ6WTPz
2Hb6bqg2/Sd4+Ri+Ok2bczXwc4EkGGgzmqWJfDLUZXh7ahfvEafmJY5e+9jwN6uYouGZDsiCd46D
VJW/OcQHqFa+xnYDGuE7U0ONGvHDYvkaex1bkxLt9oY1oLb16zhvXeFgZreqnietuqGI61lVQNep
YCCw26POWpqO9sqRWkuLj9mBsr8LpjL6h9y/P7h9Hk729oiQcDKLTpCdWz/7ogfHdDNcmCpPTbgV
KtGX5/tnCFMr7CbsrW8A1MjJ50/MCpBkaoN25oLVB4NsrPseMueJyIWYr2pijc5cplFEj09d4l4A
7ttp5b2kdhjDyqDen3jHpVLQ5E3fa63A9WUgjvjmlu6QDvMU+CFRfqGShCiqd+e7dZuUN5vAcoNR
jRzL98WR4lgEltNizgAodPWLSv2LcQw8xPh8U0KXyBy7mXFovZZGdTwsVNvi2tkPCi2ePzLBihw2
RGI1Oouv1VvyeY29b8OyMvRKXb1irihmtQklUQuJpHHt/IGiLje0SywAt7rpKSRlEHbMX0eCWmb2
7tIX4LrnLEiiA2dJv8kNMRVOFZJvBPzdY+6e9wo6ml1pBxWglMeqLLtvEm5EUi19eziTncTZbopK
sbXOFLTfFZTIU5p02ZB8GxrBjFR3xFYo8ltvXxRAGxX75rzPavvozmZ1R4s7sMF/YKy2FuvkJRiV
4BsjeZwz3B/H63Y62BLZcaD8VYhf9ponRqa0HkSPlmFQD807Rg5KC/QEH7ohh2/ARMLJdSbKlgtZ
AdOpIEjEUkoeB6wU/T88H6W2/zJDHorab4KaUXO7WqmSu/PCdvJZf7wP73yjj35gG6IkJXb7LvfG
lZNIAlLinPFPCKOLdXBIiRlCCBEB3cMS2F2Ff9jb+p021Qbljkeu5NMMppx8aTZgfIROmEK4zEZZ
OatQkBnHjjRZwhNSSfZZ6QDqpGRATHMycyggSu0qoC6me5AfU2BbuffTpSwl/SuuJwSu4I/whgRS
lTPKgs/Z3lGXZyIXl7Sga5wxwqejIS+YJnEGRujmgeJ0K/okx2kXolWT/XI/oo4dLqDxEzwjyTnR
ERq4lsc8DjlmYQ0vPROoSKfsv8xKslQTuuxbOHLJ+PCvCkP9jmk+4FDSg/xL7zCFCC2tdk2aKd1e
okSPXaS3JKiNDF/RHVQ6Ya1Og4SEsrsQxx4FmVMB2oiTx38UuNC9oS+1f1+RrKG14s0lsl4ex4yB
v1OXXGdcI9sliheh7+nhgF2Cpx7XkohaiKCPBi5GSdmP140LC24X6j0cY4ktk1gxEjU2vNw39gVS
j02EnR0Gcq4TrA8bsD8k5iwZnlcYFOMioZgdSBhblzCPS/mFG5xGH7JQZBDKNMRxavnO8kQNzeIl
KVqAexF8JYD1dp9pmk3Bie21PM6D5j5ByWUuQ3Bbq78hX6pzo4vb+gpUr3UPk5SOFHVOzFpYTNup
WGWWWZTJcInI/6evcsG0LHtDGxmpoVHrljKV6A9goTHo41/JAc+pedkZLhwkbSyU93bdn2i9ya9U
4m96sIn5TpcHDLzhe8ydzuimK0glsZ0ZXS7rL8BAtD44eOnaSSVsqqx0QXOATD5isZajvQyIQcsS
7wZy//XRsscdBub05IFEW33jk9op3TAT2B63wrK7GcIBtzMFrU4YuX562LcRBwsirjF6Xd4kTf/S
PZolBIHaC3VCzHSYPsVEeutWoY+dUoI7ZkF83UYmqbLa/SR2n/erxkaKiDJ/OotvigrSA9HH+IKH
q3X1PZO7vq+4vv7ZU/mNJORV5QAkJYjHtJiMxM/hVPPJiCuv4Skhzzbw4o7ArQ7Xp139BF4UUnv3
3JIM5qmiKCVLNaIIKI7TZAhN2PSJeldnLCIWoKHu/YW3znP5Yp8jesgunFYQMoJ002H9Do/jEYi5
W1NGKje1I9LJVkPpKUfhcIONA0LYvblhJayQxbgG83wz+l00P60V16i6qNnWyUhkXt4WCAnSlzH9
z/0bzNYf4CS2/1FKIpd1sEc1UeZ+AoNVcv8xCC7lWPcZyrTUE58tix5rjB5RTcfc98MGzZMWdrPF
4M474uZDS9TsNfp2nM7wKEAJUuzsPcfXDgY4x2JjBHRUu3ZWyUHtwcFO2RnCJ2ykmgPNNxkfrSwd
mFiDm1E2hlqzx9uumGFSlwddqarma3/Rh2dPlX11IaMpOOhJ2PnQbUbqCXzy+XlR5oZs6adfOh0N
2F1GvPx7FmZwVX2uyTQSB/T5t7WebTM5Y4fNsKK9kfRmbZ0mJ1r3ULUrrw77QEpIv0RUFS7qd25h
/i97MsKDtdbTbYHvXawIM9wi1N0xNGrNR+zDCEv/aOY8xm+KCydYBGpGSxApod74tAQwc+CCnt/X
eR4NTGnVO7u7H2mJKCaQbNGmdgyzR6VLpXaJoMnRLqBqaCbufBXgK+Yc/ZAII6LdUYVpQudNXXYx
PM4VH17fDz8INOKqjcjmZaw5nNua5H1qGPeOsgctNvCt87KeHiJH8J4X1gtwJiZVG8VMywzGaXSr
TUNIz+z4jboB9nsTz83fjvVg7BsfrNud3HnJ8VjxBQgRKNoJVh3hpzU4xa4gjR+96PdfkrXawMXb
BKl2yonO07ejB6ZZulgvl7/escVIzxLTuEUiI8ytvPKgDNUvF4t2Z091shC7tA/u0BIHskpFXGAM
deUiByRuUtL3hOBjJXbqrd1Ie8RiBgN4NuYG3wOTrd/ffV3bvfjs6X700LfhlfU3rrR1E3mI1eMj
qvA++6Sg3UuZ+0kt13NxZIjDCd5XpD8I2vVXsX0ctMzRCGXmY+ltPHAYTb+931Yol6gw71Wn8F8Y
oKRMv1Q5Q37nHHyketYh7YaP3LWCcIZRgQfxVU4O6zthJswKy8OfQpIvhr5bJUEM5UdMqR4gxHnx
nAWo2JcsyXdkwtygmpsdOALH635QA1taTErzq0AdvJC+B4HK+DF2GqHDhufxDymk/zQdKL5LZHGK
Xk1yNRgFGeQmc7Fg7ilsZJumEl+8+6D20LiN3uGQIlwzC5cfqeZ+QRg8zOV7zIOVq+FDmlsKSO5P
BBdxrHpHkieeu7AEaQu53SdaTppDkaKEoVddxCp25QKeh/FPmkrGfFLJElNP57ih59s6w51DoPSZ
zC/IPYwk2SxripJfHMj/B2MNlrVBzR2lLrx8ijuYEK2aOpfpR/smGXDu6lbMJan30EWX98F7PTFX
Iy6w17gJ5qoQnyXlpR4CqxF9SPkW9P3phaU7SYa7s1tonosCV1ixA9DJQxeJxM9K5appkjmZ+znx
5p5iIprg+FdYKl/WV4YWRhZVnOhTl8L81QpbRRXh9J/Df9aQFzc7358trOm6GUeirpwesJ04cT9o
mN8gfGR1hz82k1NQUwRSktEfaINiky+lGUd88O3ELAEs9xJoUYB6ZJ90zsJo3umgGmW3Eo7hh+y+
GtrEDv7nniEBcifwtoiCykFnsyRmZbxOh9d+QTDQ8aVr0cWlkfbRPyQRBQafujs299pAmVjiBV7k
Ra8QpgatuejHC6He/Wh2NssLrgQqs7TKVTGGr+sPTAhvwI3YoXS1qoR5h0qxdkcXshhTcy67QqIu
vuRZ4WywsOleTIXub0ulLIffyJ6m2ZECKnk5YmiEgwcYgBcmWR0o+bMArXAJi6LbNt9BzJ7kbRQ3
YS7xiLEu9ZC68CuMn4vYHuqjTDgaRkpiq6MVB2u69F0ASJxBzjI9sW/3XBYcpyWf9qwOxT3fuNjr
y4t8KpSX4t50jthvR38/HsnUHGNfx3zw+t29xfA4eX2tEbbahsAeI3dfzLrGAlaZLNgrGSSzWxlR
kYR+0F4jVe0R1RpF9bhyLrpfjHN17ddHoNpWwe5AhZ65/nrjcvY4jY7++O47r5KRhGFDchLY67L5
ajyrr21oEsigUcYIn+vA+CUlsgU2n3jb2wQRvPPLoLMpbJmNDKLh0PCcj05oHSR2C6o47wzjzp1n
/kiBhknjsLBngrBp40wFJ1Ph7Y0US47wcBiG3TzWH62TRKXPVL260if4FpaCFEdxWCZxKYdh2UI6
xUbXgKSFRtCc2aeVs3DpXBBZhdFJrYhESrA8BTmzITjpVDFivrh7Q6zKmT2+Y1HPutj/vx16MPRG
/5ds/M6eowKw4Hw39B4xir4lA0lZdYQHIF+LFy/f77hfBOP6fM6i9E8TqFIhSFy2XXH3Ivq/LyVL
YxxqAFnwj4bM6iMKwsy4gfL4zQ0XvmePyFJmw1kqFdpfMC8LAD7wKFFA/0AN+j2ud33v1nhLjkbU
GNjbXuebv07tBroZz4+q7ovgBPmEi11NAWq3U4wFQb2fqn32SGMJ/QSjUvLz8S6EZdhythaJ1ijm
9R5QEZ2+sV6OPD42lpJFQwx2jpl/BgQoCVXxSZqWyXFIubU5BnXTlQcaI59UbWlpP1W4vWEq7fkb
DfBgbdbIbh99DboDG0bTVBLaS41U7LJ2xoUJUW/b8e36ljS3GpVA/dYwZE/6xqRug1tl79jQz/wg
B9lj99xVL4xQcjM/QZjuwTKvyRPHjhuhBptkKOqEBEXzeJmW2N3GWYVSS6YG6642uqRCHQ6Mnc8F
Mm6Zel29vRRyTKMDxk/uD2Z2RDEwSlXdINUd83vXWsTbsBv3pX4NZA81OLa7+jxTT1iyvVY5dDNX
lF6tnkcavya2aIYKxEZd/bBO1mP0nbL8u5O2QMeobmkkRhaUyvFH3BV1PEqJHN9RiGFDs6pEUujT
b7H94FWAbPRjXi4+J7a1g8JhuIZ5utqeDuk01bzLbkSUwhmPE+NunKDi4LptD0kd1GWln+56DEDc
ZZNpRiJ2kEeamoPqWlUxBxoxM6DLPlj4Q4TAWm943I003KgHGzIdz/TVxCqvhHchCj5UdxUaGdlo
OXqVRNmj1ouepikD25G/DqnGRoses+7mdbGsoVbi+d16LwI92VhhYOc8VX16y07Ax188MGXxug8G
UhQ6eRF0GeEo8s/KsEoCrJ1azhVJdAELCWOVsiNWWpVdEaSXYkKtVLBwpqHI+Cj8WH2S4UbUtL3F
+FMTK3pVqUGJX1Qr0TTV50D1xpBLnNR2gn34KDje2RDVYvguuV+gFlz1gHsKC0kmHWfjteM5fQKP
xCT5RuoKg8FyWmw35OJbNbxt55TX3Igbw7/0DmH74EjYAGhvKRb6CAPXPZvE4qNUoWM3KRAO0Sy9
+1qsZuywrX+iRpVSBjUx759sFqMkYcv5QoeaGGtNmmQBOW8Pm4VMbY2vkPnX/J+OkAkbNLRVG80M
7lOhGGiuGoH2qbLcaXurB/MIo0o5qvTA/08ily2oxUPzcnG6carBa0QtVysb+W7MdEjPgj4RbXh6
lCjl1EtRR37Gd33paDz1MmgaYiEdV9osZE9OQg2jrxzf15xgQY7nrg1L+QdjkA5ar1oFXOl87Y7/
PX1oX0cWPn7OfkGrkr6XdY1CwH6BOC6Fxtc7Qy9Vn1kYMelUj6BxGtPzPoxAdeF6GZ+L8EuUCXr6
Ns1ox7jAFOtnvdVy0WeBTEINLLi4SznI1XjKDJBoWr4fTcXJ5zrN3tiLD7MSQpjKhDFodK9cZ1zE
D54Cym5wMiXTyhNMZzr329N7VbmS13Il/Bxw+Ec0pgVxMwSNzEwRvcRANfIRYyX8KwbxrbM3owe2
jqZ3AZOMghmSPAYzo+IBXCR95X/w/Nsq9gs48pY+2m1DmHouyr7UXwlaeAHCR41qs4lVy8isGYmj
UF2MAP2dPzFh3NtIIQvo0kkSd/U4StqsViNKNT3j1t41fX5fZFH5qqpyUDijFbDx9j/ZeMyL57L1
IBesUZ1Wh5IFiMdK2ZBCMGWckhcftOp1nbYO8Xzyrw6BRlNT6M9AdMMg6yZJ++3lIfHT8kdZlmDf
rK+ux/cdVoHg2wb4dWt38EzTpqptmONxqY44717LAFpWCQiyvWKnpbrEXowUq2ZUl4qyby5oQRTM
3ggXlztyCcHbIfZHTqNGWeXZvQ6YXzwUnkmlVfi0pzCFVXHIeuB6vT7sbGq9DyGmMzz/EbOjLS4a
1JUUfJdst/7tjxhpz3riFeH49XclWYcMo5nwWmTHst2hoJ0jgv8SvYi2f2eaCIgrnE06dcADHvJ+
XveKUzEs09m8HyZ/joASCuy5xd0vz4wWk+jrHkn0zJwQLjCtB2NzZwC6jgxZ8VGrELR0tQGMJ5BA
TuHZZzDCPZ46teVfkFPm9e7ZYvRksRkWIrOm8pkfZ0QOe2ANF/1/dOKwcoqCEIP2cQ2qWfJagl7k
BW84rpFQO1hDLJKVm3gYed4inDq37ehr8bBAuJq7gIWCN0vO0F2IHfTiUce/83YxD6bhNQfKopln
h6bbOGiS2GjB1tpHNt6n2PtF+AlUIN0qs5uXV1NHSrs4x6WZphhD/GiWBBA3TYCX2pyKuBaddUHz
zYwugX3+YzLekpWlb57Zyoq5JkMwtI+IiRBfejL3tF2G8MvkA7OTECT2ByOTqXjpu8T8Y+YGrN1G
pmb2R2lo5Vb4N97w0Z6/JuKXlmG2VFqDgbxZcYuhZon86cOUyDkbb+O0/jIcwz1As0TyvxDRE4E8
A6nYAfjM7TrHj9N8VSuvgES3FcEOp9bGagGyVEsxrJylBQXcXOXaCs1ux42ADv4gjLpp14IzXd49
mskOtGu4Zyuy1dX2rkCR40kZP6exXGeEbh4dhLy3tzcOESwM8TYe3fgILN4ZbWuSktVaCWb1ozML
cARlJzjldxXBn+a10f85MW1+IjbD7b1OUcmkF7LbtqP0DAy/K3JNGYxCQMmXOJRrE/Rw1nPMNvpd
23JFEwFc2rQd7Y00bWRYKlauBZC3Bl/PjhJ0ZgLnRTVs7MrFdma0MipuODeRoYCNw4a4Avelb1tF
t7EBiPutti0mssVMw6Qd4oRzBwxjItbIbsfV4TIMnFr5Ja/z/yIjaxoi02u+YEppkAPXOGg8dwyR
XaR9bxUDD/piy0VpG5b+iJ/QDXIGYw7O7xNbYYUPLzVNynZCQQlr0vzw09Jr9LBXPF8WHx1joTGW
DeN6kd2yoDQpBCIsPe08+twx9XjpioZQvrnG+h0Ertnf6kx60H2jI5N7bMZCB5jb36R5cj6/WRus
l4l0GuI4ZGhVPJYQpJeUWKjmMZM2tvtScHZgo4nkQUtzkGl5Ub8au/o6hqcnQ/EFkg3jPFXkSJAV
F3kDrGdkdDSx0tgcZt0Zr6Z2/2jWQ/R4HOWW+CnJ6O2GnBWEI79SBR87wwRpFfagAGhl9f63iafF
VsAr7Idd6cu6t/mdW4J7/0ZP2GUivkcB9MX76ZrOi3IKzOnEYrwCB1/FPp0M8AX0OKhpkl52L+P4
wKeWJrP/2P4CkQ/rlgtrYsT7ez9Aw5vN0IhHaudrd7a34NxmEKx1Uz4EPDsxZqWtpinIP6tGjzPE
frehxYr2Syy9siHxn0tgyBg3+0tGqdpDg2erW+MMJwaim09Hp+K9SJCc211rzTOjmkmOdyeLZTPn
Mb3q5fM6g5+khvm7ydfRtC26iL4QS8lKO99bNXTtcgm+grA6XjY0oJuolB3m/lJbWW/iRIxNMdQ3
pRpgTSjuM0iI7ZeLQxm3aSC049027EHa+K89ncanV6/mMlhkvzsfbBQO2Ip8OSYSkI+biU/yWyGB
8sQZJeipkfzOwfWbad56oMIT5LvTfl5juyNowQu4+GJboVkXpecPcXZ0y6+ELdm4XHINoPzxHWUg
ywSqf0GQa+KM4UWXmFXZxMaUXOV5fC2u4kAkB583pw8jI+EmZnnNoM90yOow4do6cNv+mGa2VTq8
h/KvLZ55nwle2LmdDi0lwDWrBaPI1vGiGrrgXAms77f2eSEN0PvUcxhF23HbombFCBABcxBr5Z6j
bi5EkoGJVv0/rkTkZ2CTrearMiwrXS7Spq75jV9at7iYu2UU1647U6GfvXJIqIb8IeiISzzI2JFE
cZ9O1JqBCUznhlimk5lUvPJT3jtP2t5rr5IgF/K0+qQMrz4IDtRSCv+u790sJWJNppvRhfYXLSyg
xW+88GhW14+EoOGxJw1V6kSgKZsfs2TVY1AtTUR0POxnbpuWR5xtj+Yqyz+GSmYn+nm6NrCfo0Wj
oN8kpbG9RtUjGjKuG86g5yIIe75r5XSj/Jr7Q5XgAk07jU/q8jgi3CU0gOVUv9fZ13JVkByXPk86
8JICIf+PnZMlGI6yV7b/aXUqicLWscrFt57HCiamZHSVAV9OHymtcOdhI0HAUv5hd9Hb0aCFoKQC
Y37Fg+jZ6/ZzKcz3y7tIUlvyc3NN9Us0z8c2ofL9RMkfnxjssif1j8HzvrKLGu4T7RQNDgCMx6Cu
SWSzNfYvvi8X5fEqiCEzBkpbj+HzkTDsZDZTDPzALSgzERbqmfl7OPYtGm+wktIHHe9UcN48CbTs
LyH0MQk+NbMbVObfjuz03zTZXkFgxxRfSz9jkHFcPBZjs8QcT9IEg0xI1pMQzgQY03jgbG2ddXES
wx1StDSg5jl/Hx30u3AZFf2CT4yxYB5E47u4ghKoYtw6Tr11+N1yFomVSqdGipa16cPjt7ppNGLn
U6Qh+s6afH38Opr2EzSYdzLR2C/c0734q/nJ/3DRuW7rhN67+4T2aR1ExQNYTlUTX1b/9rJpb6+K
N4ZSTpGTgJ+uQdx3nN+IZL69UcYF4lj3cPfoEJ6viHqx+HmA2qnBmivQO6HgwAfBqZNJOEgvcFRw
LLioWuyfCkNlr5jOB8H1Kjr2cfRqI4ZVHkO7bcTddRcNOCzy0Yjk3x3EShtaU31w4P5ldhs64OZm
HSxiKyh1IGleNh/AWAKyDFe01excYvOEOQmwjUR8V5Xhvyu6RXBpwiedaqO7XOlsRUf++MKKpAhg
pv8A5v8DkoRRhiLSaMP+KN2aNCj5klgpV7PLDoLWAIy7VEejUY1VSRo3CqodNkDt5Uaa/Wc6cbCa
2v4cPQYTAAWWrXdYYV2TF4eeMaOZboBigdq5Xgtk5QS28C6RZ44VFindbEbzB8zn7QRRHWsCzQBr
nVJXPS/ZJ0CHwHhkWdMmLSp1huNx6XF8siY9kOOLqRs9YDBnfDBGsrgY29MAN+IGBXw88xd6mu3V
NJe7n2ZLlBS0giL/qyOTMxJ48B9iS42xLSNni8QZM/i6IDSVamDUfbYIk4tYSxphwR9xjG4OImkI
mCp+Y6zgi7Xtxov70wu+7vY2h5MXq0KuJmrovTzhlGOKk9VbkvQVU28YmNMwLBhydih2c1KCNmk0
nCjF/HGIByGDZ07i+KyK7aT8Oxlj3Xn1PLrk0sSIyCPmhDyhZ31uhZYsq4Axl99TpEx1ljQeyPZN
7jCR6TabuyoPr4iRjrxo14yif01legKqWfjcYrUEdEUhS50zGhRi1iJHIIRTFkhaXsqE6fIq4Y61
zlQxlDKLAW5DoI/dk/imli1GjKPvtxd25+kslOzjRu+WaER+1Tj5bLJojIQVKmicXvrNap4Gkj3F
oBGlLyXu8lxpuILBcJCpFGVwIibqjLbcxGN+c0ipnk+NnCYLHHlmiS7Ef44MPMNVKvGeDnu0UNP5
Q774T2P2mYU9709cXygtPElhvNYBqJjuF3+kkK4lJIT9TkmwfOS0/S2kQzxm8ra7ApKOZ4XXNdrS
Ke9xu1QNjMa2la+IHzjUoFvXQczdxnT3nwat4wCvPXiT8emer7iiX/viq0+OlKzy60nL2Q+HSRuz
Z0AVFcjKuV3S70vY9Y3Ev2FbobCWo8az895DWt1OSYEgVxVUz/rAqSI2pHrlYsmBAdT48ggegYYu
WbdKOrI6WQoImE55nbqTU1ev9fgoZGkgJTgHTScjI/6yokJET2SWyxPnefcIasNZIHUsTqcdgw10
FNDNmg8Z+Z9qxrqJXHYKCAFqw7qTGPSeCGVKzlCnPNTboDymaTHd0ev3JXNLppmAwg49GhP/TVjG
kOhfs771FX8Cxbo7IoK3OaWBfcoompFoUhQf5m1InRTPwdJTdTQPQn/vx0c94x7g7Hj+2Sryvq/A
TDtrWa/NFEyuQZNsvan1TDvRTW+/F1dp3Vkcdx4Z9As+PeF2tnsF10KtpCptqw6/2yHBQJojEeV3
3qJcynS4ZtdLLca1n6ZACgkIAbOq5cciFNDvIwNhK2ZcTW3liKG/Y+Yc02mYV0GDRaEunu+GsARr
fjHSxq8yHbCqGSh5amS4ZUkKCdhZlt6WiNGyjeF5RtXM8g0olYqFMQgNr+Z3FP2U0v+XvNHYLT0O
fkO9qamHX0msKPQR9ysNsLkak7qSO/4a5r0pTqXt670hAzbOKwztlBa4PC6oc9NjveIQWQKrnbEk
mgFAi/9hXHO08o2iwaP8iesUmViTm3OkHmLiqMnDJ+L0ZtL7crQ5H4hlXlg5FPg8nzkcJBBKYTOe
QlM25jhRm18v3YVcUWE2gup5gwbvnkpILyJ4wb2VVKESiJ3IrRhRk4ogQ14A2gmUwZZ3VlWiQ3oA
EBqt1rCj78fhn+7a7/HZbI2tlENPw2fgqo/TkBbZd3EGeag9IMLonCLdPgNvRDk03rXNafjQEwGi
dYZ13ZOY65BTZJhKOEIoih4Hv0+I8imo4qeapTWZ5LljD/29iL8oTmSgoNttlO9ft7dr3+FB3zOz
wMjgnkc67zpToFVs1h8o4YjMPaQB2aYNgHFRpFpt4u1VL7MsDjUu6h8Lpy+D7/pbq0Fdf/CbJLcp
dcFaFMOz4YpI85TUDUTi9oU9drX5EqvQFStcm003cdhF2A0ajY8PCv5G60v8eqP6V+SQEcTsGDhq
pEg3cDnmbKY7vet6Ex6Ojp3DG8evoTKyTZcLpdetmUZPZ6ccbGT4LHL1YbQhA6NYFVugBfinZuBX
iQELMVR7JvxPLQM5tKFiFGnx3z631nzdKmrk1YI6nMhb9GetCWIl/m31FLcNfGxEJl4WHoNhiFqS
2Jj586h+ACR8SrUisYClqddC4fV34S0Dw0bSKfH474heqgIAd5f/BtB/oq5BXVMfdFVpdxoo9rTW
Ag8FuhLaWErJhbVVgbdU+XU4OxGWZy1yr32abI6Co3Sr8fEYsbN6uRet4Bu3Vh6UOsXtSR3K8Bkt
2r7s5wyiTo38kUFAolLwdmyfxs/RBqHDqwn51BPHZl8dj+SQAU0Hm0AQ3W6/TGVE4K58pa9HlQQY
27TZ+fHpBRtYGMAQn5eO/A/pCNQN8G4zBhcN81GPUtA8yazWft4pgf4N0BqeQ0+Z0SYwOEussc4C
qJNUvlZ/LjoRsjdKIjaDNizbptS4Xr1hIrk+xt0PdDPWjULEnmaMc9hP3Ki7RImhqCykEuVEJy/0
XHhT9NZvB1BHGdaXZvg5AaicnCXqvqy0M64AVRxuzw4dLtug8X71dOyJ2dxDQn0bhkPmlUUnqIZs
uxN9y6czVfIC9MXmt1ikuVa/eueHOKgHgY/XQltxzxMKhx4J8AuvZzO91IvbTk9Wrdz1cgNIUj7R
KZgIGT7JMBD0g5v3m7pm1TW1u0nNoFRCXaDxhsJhMAatrqm4cYEOvPilHA8E3CIHePHyRr6GHonb
ESYJ9Rlyk0YkWwSOgBzrXpOyaKFj5ZeJdnYmmPkErnNJF4mq/WQJu6e6EFrQn9RBjrDqptwu929L
dmF21gjismBo7nV5hKF50X39Dpt2zAgQJQuOKJG1Spfhhnp9BoOJyYsjPj62Ll82jJRSPhygmBHf
tPzvjLqF1geVDx2GxATRLo7OHY+VL/GdjLwbMDTGkH0NwZYmdc1LT9ah87h++QR7P450tOq40fsZ
+Ogzj/HR/+ozL3Ta5Vl1jLl4hkpz5VRL9yps4sOZ+kRuucZIjCdGm7nmKlwKgEh/hov7xekFj5TN
IX4V1x7Pgy9EIMPuoGZoUsa0Hads+2K03+SftgdwvpR+GoUsfw/8MamZMQiu28IJZxe3ZbcyOt4x
msTFSvj4qc2ndWTmMbo/VSxpTGeKpOXc+9+AGSy+q4C0YJhZPy6QVjq/8bz95CjAZNq5KrdBl3fF
oTL4lBCc/1pp6VbFwV0W3w4e/pNPClyXwejPcc09zpN15zNEd+Ud1uFm3R+OpM8Tco6KLD+dcFHL
8k8P0dDZ7NZfNVAB3dYaTo2a2nEeRITgJALPVlBkmLALTHaPdPk+3oKN9bPBJFGNJ5XqVza6hjVm
Tl18+L1yl1O2wEAUSnpDuTz73jVqLlpojuAHJJ85fbW5fbW7VPbO9fT4HZsV+FBztZLYXNFC/mYQ
zvv7pCw2qmNOn+us2IkW6zYQLn9jnHDOhOCbu1U37ogx+q98KhGXVla5FSQ6C4fPT1EhZUuaj3SE
lRCPMEtpVAnFIa2PwEbH0H2tLZBePVrakKJC6udusph6y2w+5lu5Abt2WopWpWmNG9KuYPqZwu6C
p7Qe6jq+7XYiZqezoL3v0ma5C2/DcMSqafjb8dlfN8XAWRFIfU6v11KO9vfyWlLGb2mA8txC+ROp
zXkW+yCtjUD9o/pOKPPuGTIXrhPyipdB3G43l/JWW8tqX7uulh0Ys03/Xt8RllST/pcTB0fokr4g
2Y5uBRUkxny5ljH3esdImEsXnj3QAKy/gpQIWt5W7JbJGyfgRxRypiiTkhE+Iql1TOe6msh/jXtX
LM9GLPHxb7HHLHCLY3DBT2knOIWlpQ2ThT6m8fsyaAYCMCNfNbQCM/nTxPViSF296sc6zCpbeMZ6
BbhpOQfJNoLKO6GoYzrIKI9QYTMouGIU0bXGPoUF5dkaXrCx8Gx/2qInwuAq7iyawA3sAzrXtiRn
hbJMSvZ2HS3LDfTraBL9QSM5Ml6KYkehNi7N4cemR9jmqnaAaxOBiZZ3V3EBUgphoXuHUcM/SV9M
o6MFGzANiVhYExoCyqHsnfQgsTUN1Nbzt5GdlYq5QChUiUvcZ+XC8r5lUHaWdZ85WKAeDovC5/3V
9oGIVRp1L1vh1oo6+3ShJ3THSOOrWikbCek6G0hkYE2n6Apo97tX4j75FGwpS2WCN8UUPVPNRhDf
8G/dlUNpX+rpE0QRdp4HFitMY8SckBK2d9rjtiGHdZvFe1HZwmHxhQkMZ7Vr46i0aWqlkRDlvc6/
XUxUhNdv7GJ9enjU9ry5jST3J2/ptVYXvvtlmlKMfXaMNVUhLkNUqtwFsidlTerywFhLDNyuZoeQ
GQjw58I4ZhAU2Hy8d+JBcfJbQJhSwV32TKumWIDeIBMnAkCz8K2jrb4qYm8a2mMekb95fiaqgQVz
AQy+/XKEUbs3BC4tinkaWTj1AasobIA+J1b4LxD1qJCW174d5jXTgJiPdtq6rskxkzeXBConcaGq
BzaJO7fm48setRSAwbLrL97++xGf61ZsqTfiTU/S37AllXaCm9DS843YsBzqjNOs7rM8Tv8YiluC
C7aCtB90d1qfQr/TNTWVPOSJNZhLTmJMJT0vpr84xG17aUaa9TJN9FHdHR81YKb2vA4M7u/NDA0+
6DoIyHiiOGesridU6UJUJwsoPTENdQu6NTHkLuEl+R67FJgmDn8tVeet8q1jDgVp4gHleejshhd1
yJsGrES5/hYuBxwdqZZSysspemALCZm7rOPp4KXLsvJf4cwjnut+Exw5N6p6jB6hAlogLU72ILSO
aS0aLx5kAnqQMAgl3jsTeASsI8WDH5SawWu9XBZlHFPBAjJLFWQOPPIgFAe2NdgFKzC+YqlvU9TO
CGZZah6qvjUM7sx1QsUMphKiKJ6Rg1t6KyOUX+4zukITLiAjnchX1yDz5kYiAoNisb895qi3No/0
LYzmcIm6/XLmqc+cSim4Hdd6xQPUyie5ZOqWW5LmM3htlNuLHJPR3Q+EI4FN0urKZXTYcSkOPrPD
f0XSakYdKdsBAo5AMETTS9BEXbZYpIFk3aFQqbQTDWbV2yAUiL6D0bC3O5JvtoHnjzaO2+BgnCnD
WgC1I8J3sj6Vr1oOK6q1wXVtWrYTMPnoMjgXtRD+qsC/UoqXaKf056YHSq7R3iSrFdE2E2X3gzVi
07LXgELx2rACv+FW9Gfs20hRxVGpDURjkEcCzYVSxBq/WwLeI4jFtz86AThvxoglcO20ry4bz0uA
VZB5PbFxyxx7cX75JnMSWBxrIgjaq6cCFAU8isvKHua8/g8fNJTqEERL8nqUQqRNAoK+b5culcyZ
3XBlBS2aygGo2Ctnr1UVjvO8+MhzsYTrG2G7+E1Rcpixw/+l1MlGq7/7mCNEumLdHk9iVcVr7E0j
r3vidy4IwAaPSClxsGTGQIOkbbi4NVYjSlwkmnrXKUeZfe4hIxqBBj8+WiJligOXNA+3ltvZBRAi
pwEqPa+7y3Z75Yxyf7F3yMcaXefNU9xKWbGWAyrV5aAziBYv//9QSdzL0aNl3IS22Zt0akR3WxUd
/l62ikTyNKRWg2i5BtXhk+yAHfhwFomv7rf7Fj+5xlzkzm423p+/ferFMLwqNuj8DnOvUxdZcCth
N1/m6h201o/9p9LtXdQKGRAXSol3rJaUhp8GlFKp7R1/Jyh0ND1wtqM6nxt3i7IdAnBbUp2+hoDZ
OtxlkNL/AtlB3UTKnkFgZR8e6Hr4BPW9BY57YPWMtfmgIalivgVQzwn73rPOHGUIEz5El8N7CzmD
9XQD0mgXZhus38//JY1YSJORZM1zNrpz7ze/TjYAWoxRWZcAoSc5/L0C8hWrZkaHEJB4NES0fQzW
j1E03iF5hKyFl1gzVrD70PvDGucgS4gaAR+qYnAlFmiadfMBgAQh/MOvFmlt/u6MNC54b16VpUMx
jkUBDmGjz8BvPtq0nnW3GU/MFHktvv1UdXvbk9ekCj/fkc1fCiiZ3ua5tacWvlpYPmY0tkOpPic/
izz73E3XhEcNpOpXiaBkAzic4ZavkzR82o3NlhBwuS6IkGY2Ulm0jkUJhSm1QQHitoZTaCp28M0O
OkZMS9OLmURtqloUQNIa6chjf+4xs6aiQ5bGpoZthkGOvtnY2vlQAOqNgvj2n5Q3cHg/9KmMyf/1
gh0xDLecipxgTBUoBH4OApEsEduCgIYRvEulG4kd9ksG1ciC+rlrZOd77/ZXmEIH2TCRiYp40cAK
+nHg/LglA/Dr9r8SjZarMxkz/qSbxHXN9DgqZbISxgYrQzM85qD0ig7ptQnlcG8ilaGKvx3/xNCT
pNmEt4XlabPVRqdHwGfE7KayyfnZJefDUbhTm1PuoZCapIXsQKt0egbXyNVMKT6qfMRpQJfu6NE3
9GXdf9pOLK3s4rzUcdjnnV8QpogBO78yv8GvwIUATugpI185jlC3QFulhw+IaYUE1ZE9s9sQB2m5
OImyZR90TiQXgCIX2wE5B7hXJek4Zcwqh+bteCzyWss1SCRvMIGarDJ8dV88svwD5bz72izHj7M6
BPbWvi4tib065P3CJe2O+FFNKwPfskUlXZ9n254jVe9xLFe6tIjAYR1wM8wQY6wK9AUdn+z4HDsW
S5eqHuQqTdSbj67JAoIUevKK63sYqMRP/AV4KZWPvyZAT/0XI7NwP+j4shjFSn1xGaugrdR8S9Px
Zg77d0HCsP1JnyN0w6Ly6vRK04rkruhRjyBIlVVMbRQ9RB6KU8cjAbfzaFZqFVxnOQjjvWTi0liT
67+P8xWkagYDdA24jN5iIaKFdzuA5fxZxQnEW74quFIqqoT2K+1S6ClFUsGVkuOwNR55PPNHAG/D
jd1Fc5MreAynTweVi17/lXZuDdd273sR/+x89j8aYFXVN/NvnQ9oDzmg2ygiRenf71kYurlmBTKK
JzJ0R9zRP270E+cLCADOJ8Oavyh0SNN2dC1J8cJASnFg5+rcZkfqlw6fnVT8u9jQ1OzVb0/wcm2k
dI9gX0rvgWjL07lBAITPu7XnmHs+gViNAYdSFM/vG0mKMkcvkB+zmH5LHDZZO5FTxptgiGK/hUHX
mTfUPgHkkiCdKDT6ZpZN6a/F/J1cfcqLnwiXIA7z/7rCSsUpRX1GazZ0g4HGFLzvEHLO1BhiVSrx
/8FeqQQxhDkA1PMoP5efr87a5x0u1t0PX4paSvDMyvDoyY6683L+Jo8KcwQGduGRHV2F0F7BWwUX
nqJHkdNdZRSFqkDwvtXWzlBIzd8XC8rOIbsuyi5Ed4VWUdYuUeP9LAHgO0A3k3LEu4dOSNVsgk1m
5tRxsaoY7z5eAUpdDSBSc6nojkxbiUAMrA46JBmOdqFz4zB67zm5GkJ/D/+1xPKp6vc15XXxrJhM
QZSuStIk1+ULd3xwW1NgMEKwDKvcqkxx6h1QuYQvv907HFx0LcyjTAzOE4g1z/ziAeBzLCmhad8q
SRHsljuU5Hqk1Yt0XqjyBRmJZiK9Tkvw31FcRfCXxQebgYTsglWlcmgba6Gtnjvggv31dPbimwhW
9p6jz3aW8sAiwGDDaZ7w09w3UQoJ3Ux6t60wffEHJ+scotokWG71039x0xhuVkpbTGioIabFeFTB
2nOFC3eK0EyOVOEpAai+id5gaFQX3hAnA/SCW1daTEztP8ZshiSh1MFNxQVRQFgYBR2Qet7S8ovx
VkWObfilqtxt+EI0IthFDYuxJ0TwARyDREo/0H9YPzrIf1i9Drk9JhoBFfM2tXj1nFsKHf68FX1I
jFu20cV46G/rjrJojYJFsDtkMQ2n6Nk8yu7qZFGfM7UZ1ZGGnAzJIGim5MgzKmsr+D1JJrsrQU+n
wYnXh6MWDhc94IPv/aW0cMhAwQB3pUNN+1M7wvDhyTWWANBcF65pGaKSIGkHyBRnhmUGcdeHizBJ
xmCIhVrEHDw1hBhditk6wUqRyJZZMC1kusTZLHaSuYaAGNgcpuOyzFJs1Aw76RIdM1zvDocsh/aO
2DYwWp0p6/f6X8GsDV5B8XwHIN+ub98Np/OnxIEkoB9Y2F8l76kk3X+Dr6oxjEMMpnzEI3Z/I+EO
841oZHV32pOAyJK5fj89QQ28WWOdRpSJKsyrmFyLLgc9OagwnCT1P5WX+SsG0O5OAj0PECxmtymn
3zESn8LtIP4e8VuHcKVDYUyDJU1800ttb0Rsfd/utKQpmA3MHy4utfDOdOQGrnPFXQl0Kiwaajl9
rWd4xNsrOP1dhLgrJ62wpAApjGP0x4kIimVsIn0q4MNIz0BXrrAWfYw3kac6btXQE1pdbn33ha+I
x/5upJCi5PZMJHT6PbRgady4EgXUm4uz0nMdcW79Q1QZFJjV9c4Sinxx4XqNIB4IJmPv8omzsZNs
JWHjMHOBTQRsTVtJ1UP6PIJn+GHSDcSTLA7HovIql+AJLS2uE572662ktJj4T6h+jJ0iNUd5yidG
za51xVqffeuhKjXCwbszHY72WZ//m5LRezppr/u17uBvToJAA6qqM9bR8/Rh5OR9FyjWFG0xSRMB
i8kdvH3gEAH/vpkfhqN4KHe/SJPpPMiMZE5ApH27buLQG1xyyyafzdlOIvoOmkMDKs6HGzCIhf0x
DSFBCoWFrHwoeqeEFMXPLb2lPI21Eaz6lffXVd1+UTnuobSy4JL9pwpVKsE9q94euBtpjaulquNB
iZNwWM4JmHBYm+FpSYJt0+dqcvNouEdgi81uW8hAg0LNvaUMAGJtt7feOUi4gLGmkwyDfQOreZqK
jNO+p0b9BW5W9/4hB5jKFjP8twObcb6zpxMce7cAn6XIa0ZnvgwuJvcHhaq9dwVudCygJXFU2ba4
h1DqVcJR3CSWl+/cnH2e7/EE9cjMwMX/4ZPn8I71tjit2shGhbuUM2CdqRlID4cMnJPoi0rJbyDF
3K68C7rOSEcCYpA+eOyYIzBPvVoL8IU+qvY8lLKFue8MqehCqmckWsYSESl/HSDf4kp//EI4if6L
7x481uG3q64n7SdorGBxRp0QyaFDssQiI3a9XuqPfBG8PsKJdR5SKg8IND0ObaPk3KBTiiVvZSrU
D13Uu+D7T1Gc/W0RGLZe3Q30QnMpQrmFE88tPDuTcCINqzZ7WqSXA5KWdIFtbfWi2KXrfBLMB4he
ZEzm48ufC5G2Ap8rU0Sn89U1o/rrS24uIA6Q6o2F6HScScwevnFyKUh8b6AXhTEA5W7pRhOKafj3
jj8SIDXrvW/b0Gy7OMTKxOqQnnJ0cNskKAZlUitpi/OxvVCK3oi+Lot0p+s/biuZ9Jsx+9BJUWDt
Jahs1pO1pZEQ2+2CAbdvh1douNw4CNGm5yYpPc2G5P3qY5kPlrxlOigk02hWg2sBH+VrBT4bCHCl
gO+xIOuZ4F3wNe3yhRer9I6jCQY+mfwSN5xoQo20C0ywN+99QbR9E4DsqxHVKzXthxnGi1nXc68k
zrZePPx4rMgf62iPi558khOqINzNvrxuAadYHbbz/imiNBGKs1ynvWSJA/p/uwS2KZ9MIJlyEjlj
Gs26TDh93NH6O8UZQMeIDuPIwSleJ6SjRNIAvh4licirRlDQ4hxuNfLQo5249JyeTMYmWjpurbm1
rN2XDD4goJ4vllxr29WH8Zlcw7LZm0Dkl/qtAu4b5XDTYWW0/JQzZGXwTJ0r3n81CWdBNo/8qoAS
SDluPSRzxLDOVF0+dsmfxuZ0LPXMcyRcmfqp38MfkoLKgPSEAhs2b/4fZmFfGCitlZftiwjVKmqT
owDY+tC0qv1679wjMKzcZsEF7DYD2tHA4Dt9OOhwhKiUltbJhYn/3gD4+pJnZwzJOVpFoyyBYmhw
0GZkeZTK4nQjWiU9E2oPi+AFiCR3B6eaxNLpI57K3gh/RJzyTSMoAV1x3fJ3ztQzlmdAIjJm4ol9
Z6II7JB1R6KDrr9EnGMaUb1T0mLCv3zbWGcDcJipi2WzfKyQpj343/CzqMFQWenSe5f5Fc25ZVCX
vCC8GkgehVTaJZalkIaI1auiCf2YPX2UcQ7dCD3HbbECMctabpPmveU75PQgbzitOFO51ZOhIIZb
gesBeRC5KAdijrruSw23gQBPkbgqRQE+H6bLb2gueMUsiamkFspHUgPWQy5lxeVK0oQhY6NXr0V0
Za5Jb4gSRwv0j3WcYwSRt1yGtN9TaVua8DRq6JxjQgZ80tyV4HT5B8hiujTi9ZQvpfCnvofBcmfF
MOQYOP8K4jJJcLUFGyt1dDbP8D343gj5pUM2CZ4kKt4WOE2lo+cegAlXZslMEi+GwudI/2Ru0GGL
nzW7G6CETWlSmYRo6kauIoetRDWURg8rRunzLr2VqAnKVyjvX6yRjqs+rly5JuduGy9pg0vrahFD
fWr136wOxketmeUBX38ityaZjg21C/uuLpqPJohFKj6e0oAWcxAdVPbsaL6k2qvvbyMd6k719aY6
zOo16IXPdngvE/iCV2+ILlqHEvVJ0dT3e5Zz8vboAKyXqIYnWg4jd0t/9Y9MIFiJPWaIw07iCX8o
CpUcd/ZZF8ZKPSwAMFnn4Ocp2BDdigRGe3qpoQ9PgNHoydrTj5nazL0D1WVEK08k0DoaAGEzXRqI
iCvsCNQvt7hMyy5YnK59GXABPrT4ZqO4VLbahdfC2zs8c7NdlYS4sa2zUFRP9WFAM4sOEKnY+swl
HWXMUaLDCzTE4ntHkmzDBgbAE26m8EIvmT8Vi5IVnzphO5DzrZMhHzFAKnWpMh4iABhXZqvVRby7
GErm0l3iVjlVnStdhl7P3RXle09Yqp70i2BxKiFo9BrsgmyByfHFuSsNLc/0KcO9pj4StlgYj2bj
842uAXTWIZ7BVAvBMGLHBOnrhHDuZ4Dg51tJpkgHCRMOklbcADfqO+1QQ4fbt76t1RSPx480AhYM
Oug+ANKRxnzrKT30eAcUH5NbhAywmC0o1MLEk/aW23WlFrSrFTaw2XrgRgL+W/AG9KD1HBbmE8sH
Se29Vs5UivDjXbstPVwmSp3d9R5Kj7X0DvwCjkDed4lXa19AwNm1mqLbFOnBzXpo7O1GRZ9VrQBC
l7BXRNbl4Bpv8jt7GhcSNYzzKfVf/hCRD+TW1H+QagkJQXZq42CEAZtU5/dF9A5jmx9Q80IixSyG
n5ktA+mLNZ2EU/QGX2e6MHzK6KQ2ek9lTyWHkd9xAcNVUiJnyKQZYHEOqJuN+xQkYbvyOg4O+V0d
sw7rp6wLc1XN0hCYEVTfpuNZQWOJBoxPpZUQ3QsJXOzO2vNX7/tI2TP2YYORV/TO3cQFU/0KXtR7
XyYnkozDd6Fv8Dd1Di0VHBH51l/Xz5tjCkGPS1niWLIrJEG1rJRDk24vQcYave9OZ+nGGsoWPfES
9wgNxbGhflGmylXPThLkVLtKfrYPKqyq86g5v0wf4emVLY84KPqIXHyEQXbPEDvEaO+a9dbg+wNo
2x95XRbTMr4ZKFsirwMJodeGipbc1qiZfpYFCSGzj/i8Qye4GGVj3Ybbsqau9hQoWiQUYMH3omeP
hT4aJes+qcKsnq9Dc7kudfyLTKESeNdlG0CEZUe/jfWKbnxoi8J356D/KYG0nR/1N93/RCuMLTbH
SzTPgUvW4+J9r743bXJSUAMRKFl3sZBpPgim9yJRFLvyBqdmeB6BmhHPADMjLxgJtmSCB/0lrBe1
a0ZA7i5zznDtWFm6hmNiyh57/DPsrJnuDsZZo23Z1r/aH6WZ84uJ28q7tTGHBAUNk4Jadjc7CE+q
Z3Q9R6lA0gbhj1iQblB4CottnPHt34G8aCfTUkNVBpWS8g8mvqkRVZB+WVIP3DNruZ/aKz5uSEVe
W05CMlfkeDyLRBRbLk8yEGkcbTiJQQqzXOGzC1+Gkx2caWQn3cDLx1FPZqSlUlGsXkE05C+00vMm
wccCsujY76hK8bbAdXnzqNkvI5p8zEk4yP6CqzkvXLVDZHlAwMC5nkR3AAp7y50JWY/TUg1oJh8z
Hph4o2Tyqi0UvWvbBJV2rCXMiQpPnho9tfSyM/uZE6wf2C0DLdCEpoJ3fhg76FtLHsmgwNOEDkzz
scYWKmVyAj3NUXrpWWAv9n/MtjsY8sDpcSfY2Kbof8J8Ttk5nIlUI4l0pHHKoWcdJnhgfkOpj6tY
GkuIelvc+n03H1PeJpwQNUJsbHQmavTTrqSDTU5KLMuLFIszhjBN19A8oD8orH+xdAn3WfvyZFSY
OshlkXL86ECA+P46HMwGCIYf2mKupntrmPneYY1XK1Z2Cv3ZbaIOuw3q1uhz8WOqbnm/qtkeGucI
clIiksg6zvCO+JNmkDMUYfzp3Quq09sF/fT5ZLjN4gy9VXaVNPtdToG/jlbO9XR+0Mv8Cw+UMSjy
odYPI2ensfw3R6Wi9NttrPAkdDcgusgz7P/J2c4fXci6WdhQi773qIvxHsfT1L/5g9qwuOHE+M7m
rkwvgFQXe1i84GOKju0WTRniypghBMMnPW8dbc4VzaaT+w8vLd7cQvBBYjhR0x/g0YpW68OtyhV7
PqvSDrx7KrEcGu0YT73rjbtbjeUP8zsGevCWhaHt2r/b1CfL8MBmGUDPZw65m7wTGbl/DAcoEpWN
9hPhGKlbEGT23lD5S+5bprowSK+WaHuy3F/IrmNODi3GJqsunjX1rqW/D0bjADJO1P7otlutqBej
VDX4MqK60uFb1M/n4lU8/wP0IGVs2ly+CV/wiJNcVhQ97C2nTKV4Rzfx4w5jGlMyQEp1F1Ppa40c
hS50ELKMGpYB/OjyZm1iPE7Z8UAoGamk4JFAxOitD3on5GVI64w/DIKOnZz9K/4cfD//lK9TQl6e
xyrfhHZ6s64L+CEhQY9eumWoxidTNREl/nLRdva2+sIz+QDzBJI93sy6gODs+wVCBULsBRJrkfUa
LUCX2FXMCEfsxrT2UkxODzfF8hOP5jtCreeerA3NkMqYvvIYMDxXHlOi7N2cbi2BYKIx2YP+/1yY
yCrpmiaFPlcMKcFOmTxMLMBCHbZy5XYaHkdqcOUo1czqMyDJmgKNsC8y6DjU0gr7wkO1JxfqIMBe
LQCoVFQw8FL63GCk3Hjrjs6c7msliPH0YvLVk2/0meWvtXji8fp0Nlhi5mpjJQWjsRbivbpmLurc
lu0Qlw0aCXFPbXh9QGocClunMFHBPqpNRi0BzZY6D4hhbSzmeg0/G8TDQXZ7LDN+BT50ILeL/S8b
zpZSuI57WQGQgVzRwW+TTwERDtRYD5fLMk6/6P3deqoV+x+mp0/KATup7TLsGRuGAmEJzR3iWX3g
zrGAjI2uXnLifF1phKOV9lcZLNmgAsyit07l5kVrwmNiVXwoM0BKSCDFim6TDmbB3mQINK7Ajr6d
boaogcJXxizeSqlfjVFHgI8SfC3hanve++ppaYMsbWDkpq8DRVzgeEZhtThBTHOKHAgL/Bm0zG0i
0PHznoOcjqPjucSzMzU3BTWcZEuuksz4EA4MiHhHtrloLWiUR7ttSUxnXnCZLZGG/jnvYncidm7K
ZHSOd/Cg+5ikRaOn0LnrVRTQdU4JUFZIOynAh8b4bAyFF7ePiUGtIdLCCkaUW68/VTWm3QYmv41l
Y2fAZw6wtGtRQZ5dlIm6nKX+jTuGeO8oqvMTPrD9VVSo5AQrbZrGZdbpF9kbg/aUXFA9oLLeelQG
Xr2M/3J9dF8/AwQOP/nBD8VQrzqddawbpRdQpSMGJAtkPI8YuxsxgXfIjK1kGsBZUOjzSeoJ7T5z
6lZ9D3rQnTrtrQmEdvitkJitLfIo4k0jbY+o2dWvClLWFrXpM8nFHWU61V3jHLkgXyReqbRBHXBa
8Tj7M4pT2OAwByjVdKcb/iV1mYyjGO07u8dIoLGkafsfjDOKfdYfgocSgge4JTZN1K0Sy99mVyG+
myOEcaX0h6IP4t0+C1TxUPbFqVVTiaMIaPK+gDSZW9dwe6xilEWVuP4t++ZcKQSAEr78YNsi9BwP
n0kKV/+Y17MTMTAK6XsJhx1QHXLGVDEQDcFpk2LS2far7LckFdINZwHUu8G8VtajnVrenAaPxFPq
roOxOJD5jpYBrPLzgCEWmfgrY9lJaQq1qeWEQJau9UROKmV1IwDXPua5U5r2xX8/YA8/4AqRLCIB
5YBytY+CTiSQdcsl1vpyQUPGib19lKzBdVVHK3B3Wewges3m0CZ3mTsOMLh99HsLcR6iCOfEPv1L
UBDVRIKviV48OgPW4wA6t92geHsuzP2N4ZOAx9fHhATBZu4wXIgJJZy+V1uuKV9Ps1iUkJQUU24J
T0quEYKzyMLPbRaGTaTsYlWlDPry+f/v3kkwMmZeUY48mMyQswpGsNavhuwiurtC+9Cza+ejHKTO
9Gw7rjnKGVpSFugwB92hcaCdp1Bt5b4bpoAM2+GQNLEWtbOQmIEHRVwKorjfl4b8N06skuROjbkG
WWokvrNiz2OVOS00V0oU9BybN3W+QbWqNvW7sDBB5D0gdwcd3ONCxeIBzEsg7nfwXiEpZpMsLCF+
KLXECNkoqv/zEkFs38VMfsJRScKHuapFUUoS7DLO4Nrugj6ZCkX76F/Zm8uwFtpBYuJ5biaaLiBy
M+VNi41kXg2ku0D5PcdcY0ugpoAe+AzbsHV1gfswtqTjVtekaQwc9KE/GEPdq0nErpiguH3dMxlA
aUx70FmQMa6PF6cpO7IV1QASBrfd0oB+0c3KnsA0kBQ0Fcw/v2fdjOmMkYRxxZ6NlDKWwUI+k6u9
dc83MvNsXqcsmH57A7fPU/sdd4FgVkpOt7aGdgje1wyd4woqF9bqrCUEMluxjcnYJIttf2VIbM+b
Nl8Y51dXoJoel5qx/Pa7E/IIZ/tRprrpmtEmIV6mOfGrmhss8y24TMXBNpCiT5lX2vLrZDk+yG5v
c+xwZiO9Xwp2tljvx11OG8is9okT9+3RlWVBgicwM7Rb/sZKIlr7Wnhiks3TeyoCXkoUKgU/jzfN
BQLNQhy67ddY5v9dxaOefv7oH8dUuSM5i0/RxJpYf7Q569WoxLzaXEuxHSdr6KJ3FDz3gWouE3oh
gJufTjW1yxbKdo427CDFcXLSrr7sep5I910h/rEcW35+OkBOQXH4lAx/RkfrzqaOPSr/5A5EkP97
ANNXRGewYeizRAc+8+CZe/HC5bfSgCWVPvN6Io0S0u0A5FaJ7ASOFIQukgdQaN7yJwmZc+y5ifV2
L+N20xCKWKueptZwg/ln2wGeXHQE6iuObogLSfOnt3Y5Lf1JbiaJQIjmO/jqE9Qz6NnhsLeaxtV/
HpCRW4aYY9tJnTZyvCg8EONHUbLuPRPiUqd3qJV7J+wEqBYWZ1Xw11AYwW1qEsbykDEliG1FQQaC
LjlSzESNCb9bpKRVLhe10S7t695sW9LnJIA1IkKoV5HEZrJuVUn7uM+Uz1jPbM2yw2VbhwMhRCFB
RdgGzfJSwR/dvUUyJnDe9HKBD8wOZ6uM2SBucGDgTN0Xi38mLfdzRLUHU8Cmx9QUBVaGqqLb4CYe
pLjhuHA6TOSVxTvX4e37+4lg6P8/xBmiI3C8KtuHg16w0XsbOyQBsMCjzJwtmYz+UG07oH/8xBps
B7Ga1fNy+yU2XNFliOQiPcDpsnN37UlKRkTbXy/G0THpSMqfqeyzKNmJNWbptz8B00dcg2fLGrC/
qwg7p8WuHQ1HqpkVZqgyE91JLCq4CtM4nYJpJcN1tEe2Q6bEyj6ZVGXnZJZugynVTXrINAPYFcVr
qEMaSgEgn/76xmGZxE/kcsBgnu7Kkrvq8KjAxEZJMHSF3WoYjPxBneDkGQm0qMArKe2WCb/lSiK9
NTFZXsiBFjzZrRmwnjoMo7jk2iQJRJvOariLbnvk37srjbLWgL1Bm5Jk+Bh4naBNyWUQrm012ER9
bltrcZKdyeLnaYsy3zkULj+JfIGgynRWp26OirBI7b9Tbdh3u+cOp4IgBT04+QFxff/P9vNnNUWW
1Jy6T+pxk1XkwX4KDkEMY+xbE/aZEwtnS+/+ZtPGUSmZgXTEwqVQ1DrMacA+WUTUszyqgqd05yX8
v1xTm5Gp/oXKR9+I5PNBixM1vAx3YOjQHx/Sa5LYG67ENArKytZOc0oUxUgYlf3oKP8f8RwzIC3O
xCTj/O/ihGSA5tCdYLMG8CGbMFYw26/UN0njXiXCPzZ+dsQndue0zKp4QR0TEeyO971fl3G85eV1
se5g36RdTpU9hVyf2wPXYHsCg5B9Rr9MxEjKeJsANoGKMYyxTN8dkBGRm8d+Dx/W3VQ2aIuhId15
o0WnjZkaOH0ZLtroI0qJIhDoNVwhyFol+1H8+1SmklXRFAV/bfZ8oghM95/ZTsmTt/mNRp1ecZpd
xRboQjG9VRQuKKNKVqwE/Pxbu6uqk12zoglKaaIU8PW9skiRmloW7eb84xwDj/cwCRAqa0MNlGM5
blA5ZJp5EHL5B65QGSuGe0aIXpLPHk3C8Tmrze39ttkoGX0QYzKSfAm7AQmdboct4RsM3W+Brab9
/dW3BZt48Q7ygIXzNzsovv2354CAWl86VfTjELSkgVghjMhpS9q9u7UlJyvNUx5oY/lTw8m0cITQ
DEX8w0/t3D9cqbGvuP6BOlUG1iKwto5isiv+qkEkGV1CZx2lu6i8pkS1TDUtvM1XP6uLOoiMqAoa
bHcHV+vWkrrlawPmU4CglHPyqXB9XYCb0mnDqKtLI+BEC867NIpI9Y5h3xmgrVZkDyT9gajEsWqM
/DSLyILbHe5GUc6EJlfFSxzfc0IrwPZrzr+wVs3UDouBfcBkQNkRx/CBU+TSc01LFDNYP8HhAmF9
TIYIS85LtO9Q4CXpiPFbcRqnwCaxApsabfifd5ISrYh7i6j03jL5I0xfRjDAAe9X8GtA3+2zEsJQ
i5CnqZO7yY5F9zvYqMtWoMoClvzlgFdC4dzi9Mk1++ukQ72qr7ysSSHUBNwTUJzfyh/1jjH64kE8
eEzY/xfZZLEq36C5BdCbCW6kAx6AyTr/7n2DlI77CVxTSWMcWesKp3f2hg4fhuGFerdyPXy8yWGj
AzGObV1yldyk8jttVKocWtAzu3/MjQp/94j7AZS+aMDVVUuC8D/pz/8KFmqk15pHUTDANzXfVk1P
jKMWg6bfMsM/QC70/KYh2xjF5kHtsCnFfu7iziYrntefy+40NIVrGJWO5drpeEQwRd+QOFYKI2+F
2QZUhrEfYDPkaDWp8jYb0ugPF4ZxryVYy75l4mIL495YaQFrBa9GiceByLQbhTdvG9aDRYextYBI
Lk/BQ2MRLynroV1LbCAdNPEaReOgI6P+Oox2b+sYfbnCRblViYJe31yEaZmh4b1K7U9oFNOfQPm0
o5i2se3Xe8EsxKEb56Z0qJOp+bPi7OBLkb7iDaZvim6+2zY0/omrzLLKIC7UZ5qhUbune/7ufn+G
8zdv/TUlzBZxliKV4jRpiiChrp3O+Qt+Vti7DChn3/kMTmQK8q8IC4KFBThTLD6cXjp66oAZsOTy
C6v8IPxaZTZ3qyDxIxfB1cI+qwhVN6FAfItSSOuNSWJAzo+Vk9MxQ/tnZsUubGryRX8BNf8NPwsn
4IGCMb1TopN9mra3dElWdthZokjMWO1hvCZ+1vTKHfzyzVCP3H7Z4mWbrOVUo0QmthGqRjdWhD8C
BRipNXP8ooIJUPLh6EbyK5WV7ceFPJIgYnc4d+U1FJtEtcoK5LPpQuLzWo1CeYToiSDCpS5loIwg
JGOHHojkxF0809xUeMYRJxxCkV85suZB9Jxqxgg5h7IRndMtHn0XXFWx2/Xz2z0C3yNddhE5nrUN
bwWvklVwc4cLyXYEdA+CyWxcfZTTLzpaB4macB97dJmduKqW1djJbwvzOoKmzxpoGv9Hz4XNla/5
ufzCI1h5lFUcVkzmf70u1sfIlBVFamuz0YwpqzPgKI5NNaHqKeFouNgr0NVdOqcXSwCG+UoNOh8e
xQSKvd8ROey/BOvbgErAMFXGyajTPjlNcOP6ywJPdI/b0wze24xZihEnb08/eZYKJvHaP7R6+w17
Jh5NoPNv0Q1dKD5iE41C603qWRSi0UZVQPv1egp/myyO/XvJgiUHoNdBj9SfHlHEb2owtUr/IB4/
l5qwUcD07B1zQeCv2HA2eMXJDdYYN1YfXLzDkKeLsFyKifCMz5WJtDPkqgdfkSwtcvADJsyBP0gm
6Kp8uwH8ejSwPUZHHi05a+4OqM8DW3GVpkLjsrsD9r57uB7aCPX8Fqa6NTim1UCgqBPjRESuhxJH
wANCMDdhbQ6+jMQcAXR8B9qik/YSkR0c7D0ZX8+nIUBVazwv+f/wcCXvETWWsP9X3aPA/BganObn
26OWpJEU1nRCouAMtxF0WahJADSwalchxtqqSQaY7S4Kb/n0UEWLr8MQzIrfHh2EJ7AmCVJ32Sb+
uzPrHjgwECquXzzf1mLUiv9nHvg3+uq4Poqu046LGkML8RFNcorM562vTaWTah41oMADdTxFxy0Q
F+7Fe5g6CZ1ZSv71RoFaztr9aqAWQ2LaDARO6V6+VMh2nXmoSwXxRuKQnFAagtR4rPOVwm33VxLn
JRl5QjNroESzjN7KsIm+6wb6+LlL1m2y8DhvncNY8FaOZjpdb0Vd3rtxFdSHxybc0kISDC3JEPfw
gCDBM6wg/DyN8uglqincPlrdeOaRR6h3ZOyYHV9vqRr8B16lCQLWjP0U6NETd4AlCep/DaAI7Z4r
LqthjGYJM5MieP1krIsgnPUjBSj+8X/qnKlCuTPE+zA/BE6XG3eHZ7wr91IkCFm1G/u6ft87AUfV
ZYHgpaP2/tUfRk1yDcRr0t22EfDf3C8BURaGxzk66NNKc8VfXYaWI/+eXP4BaVK1whvbONjJ1rti
aKfmydXeJdHsab3gi3aYmMJm5oe6/zZG4Bq5halBchiCyUw5yPoHOEaLKJweb3hG5I3e+02L0mmI
77ElP0/HVG1fGLM+pWfSNEZ31EhiCZG+4rE+qKflGAIVX2zAhITuA6a86hTRLiRaPMqpbbNXBXBc
G2a9zfALUWVguyFOS8OmWTbwlrqGTANh3EWgHntLIKH8yyYTpKRYdXqAiCfESvbrHD0RtVRgHIkP
VPkbhm3826+lLe3IJF6a7MKR/01N22MS+Fh8/DBmAQOzkfBRVpIdb3UdeKexWEqZtmQWeQxa/ERM
dpcLHes2xktg8ru1UjKvgc2OP6DtlGRl7iJd1K/dDr8K3DM5Q6XXv82atXhihJwFNftIwb8fJNOX
AoVzjn/fhS1u/ra5RU9Z50wUX8fTP7Gm5HDEMmUJxPGKY5ZIfPHFZZdUanV2TWrNWe94fzvWoGmH
vZtOfWw3xMxQ28uy0hWPcuDqJTJcbX60LZqcaCVQ9lkKJuzi7YxU6GiAJjlyYzkmsUAbsrCEjmf7
awNJAIlNl6jWIh+E7B6N3KYYduTb6zZhP+yiSGpRchBTdILLfYA15PYGgblFzFBMnxMtmiN+d8Xk
ZwmEr8Up1N7s25lgtecjiFdzquTB0ESQ67mizb1m/VTCixxTXhj5GNBYlxAIm0W6+rT60phZUpEg
fERaBObXxKfaWAwra6J/oGEt4Jtz0cgy4VjUYU5zuKaCwTVU+OXmQ4d5qfGxt+q2VUNJdirdJFW3
SuGppOPJzJ+gf6GWzglviBhVQsKIG5bzQNAWTjheNTMfiU0S/jruzbKI908OSKTfMy68wuGYlRmt
F1mfdYcr9tGqlApI1MTnn3rCxg459xC4xIpkAD1x0Nh9PuwHeVLwILQYngCR2rc42JhD5KtBaf9H
F0lfn1KLPDdLvED+z6AizZpmpkXqsGyD8AUlY6g0i8/6sjLR7YnAEAj5XrQOvsmQCWH4lofKZYRo
+mY3zVm3GbjBomMP0snRPUpl/aec2fBDrnNew00fm+VpPOvjVYVzsWfrCfmmsfR8IhLeAWUNmAiq
/+h2go4CLX42+9BVmVQteGsUrEGQe5LJulFdjzeuahtmUaWecs2IGagQc4TLNDkuVbiSvkKab4Iw
nN3UMsf74ZsTKvpNbIZhnvRvhd6ZpjsXrQN2eh3Iri//d02LsGUEEYymRYXCuNiODDwH5P1Rutlx
PZUKxPdMB0bwqqdgo6LYuyb5TjACgN1iGv7GeqDvOkP/wBRhZoki8JqYh3rX93kFKYA+A4zuqZtj
U3/4ll8QhTAoEoTen4pYJPjrPc0Gd1EXBOHLxfiO8vp/ub6uojFWfYVE3HWk9jGuQvpz7Q65ifQx
R/N7FgodTU8oDrRQoKhd5oCmLSzRqvTaNhVSDMpk2tRRmTr50vQ1as2l0XlmjuvxMzZINwnBaXOU
PRyg5VA+TJOQHOJXrFBx7a9bSA1xZ7fuvneowZIvcarHYYMdeD7DfvKgbcLWMyqvH4NoT8ZNq9/F
uzY396s1KUt+tRq+XQ3+u1pzlevCa/dn7QjNtNiDQUTsjOoLcmSpQsUA/ywPgf7gglQgOkPwQg2D
HlEE/TMM2DZpbUmJsC3fAQNVQtHleEkvcD4TTLYxKFGkPrOpadeCgjwjzmhlbb+N50/p+Ma8efyD
zQ4K1EEX3uEOla8RQm/FxTbqMJwGDBAAM1DyZmhtveeLrw4FVSKLAboopfNhgNiTX9jZnztVgAuR
7JRvzhkfmgtZ1uSL2HxlHCMu0GJwRfTLF/eHo7Ym8G1ef1y4UI+b/wXv8seV2DZPM7ryHqzCNCHX
q9I04y6xfV9R82D71U+psoRhBr92B7nMjkrq5jXsJazEv9qG5fVhHzf/TrtgT7Fq2rXa2AQk8cu0
4r4CN8NysN4WAuk/ZYIPOz+TxKguSZePuyON2zab6mRebpl2egDRAeMEEOHjJxgWtr4SzdRzLlkB
gMFU6MenDZlm5UStTcRRUlMBA1LAbowZKRTmaoYRvo+N3o83kxJALPT7A63TDsdKaalJVOOlDVLM
Fmx8o4EoY+WnXC6NmMeFOMIn+KgEQHPLaaoS33IL4gTDBBIZ9OFK8nKOVhpW7k6LJw27yFVgfbrf
V3M8z5jwD2gW6em6rBcKJo9V6jGhc9rE1KEWe5K2afHVymCXijBwtdqc+DonVzxikIWCmEwfbt+N
NXts1o4fE/Pj3NLYZ1YsRYR7MstYDePjN2JFGNZ2XkMpbjLf4q/9kcghDycDkOqTu439j7e2xofc
sGWKB4IRQYkUrZjMqM8yAmLO0NnDmJ9p9mpRqPsIMuPp0+1Mzxm6cwe84megsi9c+8surh5WfHhd
xYvzKlsQ1sL0rHXkhI3/Gcg7uvA7LheCyhfb7p0Kebyqo+fuxKBCiGgLNc0dlaM5BI/2gJohQKYB
1G0557teQDnLWAF/WMUb2afCj7dXOiuLB5qjXdDvTVhu+/xEebhAJJUgVTfmVRmaRziUAw/z+ExS
IJ2W6p4/1hubPdAL2fp3ClnrB06BEZxLkw9RWh5/p8T1I5IfeLPDoxnteEo1fP7ApLFYS71mFCI9
ZQjRpEGeO/juhhzZ0bPxPnxbko3fQ9+87ot1QhFSORShAbslek9pJOTkeZHZB8GOUEPj3ARtcE1M
QVmyx+kz6LBiTzgjWU4PxeYKgn52ZwlZUU2SlvQEhU3JGNPvzrrxYLwwH6IfYnXlm7XPS2LrRlfK
kTxHLN0+mnmZkl3E7cipIvWO4Qt/IEFwgBap7AD6n5WUXe6G0qI9dlrCfIKIIHekTcitWqbOiLZs
97eC0L7z+lS+uJu98VJqwrTVWohFlhigK7DpCi6cefZdrhsiHeuaue6Y6bcvoh7EMm9dgWKPmHk0
JeWfvXspCtVKFKsWQwUovYGV0vFbepO+26XGadpBZhHzo56059l4CZvTtfhTMWtvOA7vc9gGV0a9
M/+J0DfbQVuhnp/r1e85kzLAGuONaHfDMh8PhTTlCk3OABiL/7apUy7m9kD81DDJ8CdAb0UOS7E7
GwiNK8iwu8h3nVd2y1Yzd9vWEkfWngvc67BlaDdmBo1MKy6lWFJ/1eoXbFs770wysDeYB/wMJDPG
g1VfeX2mzyOtvzN/PDxN6KW0zyqtbGE4T4S9Ftd4IuH39Ago2ApuPtMgzeX3hu/j43QBNu/5+u/1
nk8ahYJG0BH/kYw5Xcejp7szcJQI+LkKlfoRlOzUTlD2AZKsRXoKWB04VzwNdBCn400LQ/B9ikZ4
RwdLZLq30FST7Nuod3kd+aIsjctXlfjJZPSfivbf058tSRMfzrhXPQVCEJyy0XodImr5B9Yw9/Fl
kvnfr15fL85gSpyx2jJ9H4jDoC6lfPN8ovwloWVKek7kUzDAzA2QWtU7+LXyqlAYMp22KUE8nFvL
ezmOmdzNwi6n2gT/QDuuBAivK487SMoUp1XeJgAB8dNxZ/zZNpcvpyyr72gpdtvTGh74n8MMOuxG
GAHgsCvDqjk74iK8TLsv692OaRR3mOrbTZgrENbZlXipwQ2TCPHoeN8pZa8YGL840Ir5C4b/Nx/3
+JnQnOPwHsZ/BDL/CQ7gDNmDb3qGGMvQjBBRIYz8XAR1YM9Yly7kylsmVoxJgLyjg+6m08xwcM9Z
mXhw4FkO33L+f8to2iwCW7meKeVPBYh6K5BKXrlR4TvixnByPWXPevuz2TmzuZcixs6zI1yKm2VM
gX471TV1B7e/UpJeBMYoxTGJZ0uBP1IlJugZBotlayX+RZhcBjqNw8BUHgM1zUA40hx0rsYsWWpo
9j3SwFCsOQ0DxwbGLYPejRfF7My/NuofCNQQdNubkipeWOhViEUkJzu2mL1yeedjQAR/i6+NwGqj
/4na+1VxQG5QGlonP1FpNkWf27W7lLTCJTdkncfRCngmJQzL0sS9vQC6mJnqGeQvsDbhQnio01P6
n+1Hpc3baIwTUWxi9XvY9T88MTI+PcvJPHUeOv/7ao2gi0VHjSW53V0i8ZB30r+oFASVpeCKklAA
aHv+8cfd9g0aYjuMlnFaKgCBMwm/0glJZk36FT8YI5OABL8VPE59yZILOvKWIIhHNJ2DM2bD/tpX
s1kJIxvVeMvCnmvZk7Np4UbiEJzQj0EKt9Dczwr7hbTORVt7eKCt6NFLewbsDJgPNc1yXkCyOB9T
A0rOJYCdb6IHUmznagcafbBFWRe2ff7NQiNFBZFNc7L06JncETB62HZ6anhY9ULdrbhqhJybtkvF
J4oC1Y3EE6jOlJv12RNmDRxYLga4+Z9GGPE/KsD+iNArta7I/aGpHOwIIYbC8JrPosTr+i2yFa1+
jy8OhN1Pbur1vSrEUAfkQ0sSINjYcwSdr6UoUlRvLgzB3lHLBr0/aSJAM3pLxjUvoJRWiC9QcHIX
KlMNrXxyla5Day7rqTPtVfqL/SbVuUfmE20M2+/Ur0/6x8bxlfqApaT+GsyJK7LZCPPJtercGAVR
34ldQY8swEP+TTdYWBl+RvCQNi08MTI6uxkBHkzkpvg6u5YxWMufB4HV/0wMlFvGJV9dJwnnSsXC
X2Ph2oXqMb6RSsu60NpHFSU4b9V31ANm7zerNIFb4q1tIlbs2FdsMJfvJU25i/gjLgndG+Hj0SVN
NSzcb5a+5LgfMSBTM0VdnM1lv2ZgMeHL3ftlhoG8QqqLHjqlDFSRi+0v9hwetVoSLrJdp+kcuFql
IwI3/FW9tQVzl5jvObCfJFRgGMH3C6CxFjuLlm8UMLF3NqtvCi6TbwldjkEc7HSBiHyMqSOIzBB0
E7dghc0dpKK9zsDsvcCqK5E5lHzMkmjnIkFYbs0TPP6strNlnOSu6lAK1q+qjFu/k1eOikhKMp42
GIQbK2qi4l2D8fc6T91lIiUoF7QtO0e+25WRi4NyBsAvhP6KWBw47OnI3u4AGTeszTcnEi8gJj88
o5fddYHbqptVwG/basW2EmPF4c9wHJ5Y+Q/l9iWJsXoIGuyAjKO9dyIqvGEKEcwue8qsGZ1uRqmp
y6gmQcfeO54XEUr+Q2O3Bd5wRRo1v6TpPARK2skmIcxA1fMrG2PZJ+SR4L9Txh76RG0sWW617wCM
/Zw4gDfmT4jPVh7O57UXvCImgENp8Q0/oeJ+237EstpdgFm1dTN8tQkSGnwTM9JJy7C/6F0WI5WC
0y39+R4P11plfT6Uwbx81pG8vEyO5IitgIZBJcHphA4Y3dmb//i/DyAHBuPna3LsobKmAxZUb1Tb
STT3GYrGgnY2EaD8w2hMdA3JV3+HE9rlepnUv3SkQxV7bwCqwk+jV/A8iZj3u1HEdXLQ9lbR/tJZ
GAL177r5O+an0w9RkLZoBMz5cn25A78QwbqznqNBdiiO+PLHNStvPCkkwLiAmKg8RZvcaW+3Vhpg
33x15GPN9VxoA3T30ZoySttPy3FNjZjcwzhAmc3er6exqpAEfgDDsA2QqdBMiERKWqIHrp7E5Ue1
wZ5opnZfEhx3pY0htmKMwgPAw/FAQ/MuYUWuvQ9s+RXUqMqX2c/9ipoIul33EVInzHgncnTEuEO4
mGV+ZsXaN/5hkY6nHe1wRTCQdOP1exehMbVShY0QxL+8TgbGr7BjaJlkeOx9RMT1C7ZSaxJfmC0g
rgFdfYwV1Fh58BJnyeeHhcKxWu5Oz39dBLZedsbFoB7hq1gVXmR4ChsgQk2kS/hUQAM7IFRaNPUN
2n2nw2wyWgZ2MdzBPmw4/ae8bLZC0jMPyh9URNjzIX6tTRBxzCcOhvLWAFUWZE4JIDTEooWjv7Df
lkGCSjqkzmkp3DxhIi4QO+vWeqUmk49E6wAw5KCPN3L/T2ysub5AhkmLWFe728HxODzfyJJ6Zx1M
nr01h6FNk1eSbNWwijgTeBzMA1oKvbs7bLzNyceoCk+TQD8q0WNDaz6CTmr1wGA6/y7LNNO41df9
hrJWMJLfz9qWlRfb/D6m0BVwy8PrsgINi5/bxPswhJToYbI/nxAyzro3sPm4GClNNXItNxhL326/
vPp9vPEIaMMXgYnt0VVP/PjPL4TiJmE2ICHhesmZC0QLhXXevYvlyUZUMF7DPI+GV91YosKjUNBV
CC+knDW3WVP+Al1JlHDvkM/y33gghPDESKTo2yNLOa0vY9HG1jfRPeN9DtrX7dIIHOIlz5SgrFOm
si21PFq0O8awM+b6XLut9oqeBPagAFZH3dHbn8HvfVH3qgJKCJLHYGB2e26KAhxCnktBfwSjdkvJ
DwTSWAe9FM7mryU7Uhos5jlygEjomVj65KL0msxC7f1QTCxu3jugzq0xpmssk2P8bn6aU/L+v3ka
FrTFxqJ43XlV3Y/M8sxhVHzznYOlNcMs8NdnOq97Z6bL07RG3GV0idJoQ+tqK1z4XBqh7fME78A7
kPvu85xqRNu1JCv+haiFnmmlu0TxeV2h2/N7I2RTFKzTtkJCRUC8jGWq2IthaXP7vnCzVoH1hekB
1VaQMLeOW+BwWLyRf6ney8GfaUA8fRqL29/q98xIe7Im2b0bFtC78Y3OAOIHP4+TDr0cl+WJbwea
75SIbbkHYsRXKckHTMyW/LRhActj67p9EZ7GI9hYRuFt9IUgafGieIVHfCQPlIM6m0jrTGi9LDbq
T5hRZzlcJl284fNcFp1+UMRn68Unx+EHamHeA3+oMCr7BHC/EU4W9WtQkurAZJfn/hLkcAlB/dVe
VrcAtt31AgSW41D8yMv4KDyqRyEvDrS8nAciDtsI1PyU4NZ8lWVMz3LeihlmfZaLiAPAeN+UdQ+k
cTal0ArD8C0TshSTCRF//oscZeiJ42XKyWMjaMPFQA+wInrELpbsihDmqdYYjHd8SetD7nkgox8/
8Nor0aPJ1p3/LZNV8JWAd6O4eza91qgctsBlsX53pnsI1xqJQQ2u0ceZ0faPpdK/ROm1vwo18w/b
EiglxyNQmEXdhJF9DDhAXGh8tXSC9axrtM5dz0zWs2QUqJm8YxPvMwDVI8RVGO4KF2J8nAQGxLtG
vhTrmxnFV4xRY2rbaEhx/bbe7vBHEwovYaU1yTJ02UysPSrDgG76898o5/rADFs+fdt/R6s4TEKl
j/yycROynvFf/VJaw31bI8XkslETb5NdcC+NUfyfAbAqfyqNs2feCXtEbpGmQshr1ZBvJwO4s/kz
zQh374n38nfmqx+xEfpgyM3qTox1lLY31bxoWsyoGw9YjYnOD5luenH5p0dTo4RfF01zbAy7Ph0G
8BG3ayozx5hH5ZFWD4KH/aQ91wlVZk4mAthL2UP7WClFDIs3A5ktXl3iqeQFttxbptDg/+RCO9on
MhPgNoKmJKscO5JCSis6plqYGDOyGM7QZshjvxyyir/tgfIp9MuXnphanCgoOPCYTLlnunCItImw
d0TiLpX6aOd5MYQ2aJUVuwdmyvRg/knjTpy3rCal/O6vUyY7qhzOgLVvV6UiM8qqIzf2iCcwgKeT
D+IAFnxwrXW6VkcJ/kB8bFuBE5ROr21Wb794cEfrQ8kbfV3bo+KUR29SBQ0+iTE+xyI6yzX1GW5d
mT2xBZZWqfie3tmhtVKBqY/Wu6CNc7eurlgXnePWc27DZAUEyMn7/UAPhJ1WkJEDF8AQNxm3XnHp
mK7z90MEIzDGwRlMDPqZauPNAhbof0RoehKZKa1anwk0nh9Iw/akAwGWRGmon/eUj4zrym+GVP8/
X0Z+EiJsag9t8AQEbUFJEO8uk/88ufxpBRJTzWdcuLVtDsUCI2Ascp66Q6O8uSV/O6nCv6I1/xjN
pcwAadj3IVzHxJlx9g0tmaqWQHeS8wgdll9Y2K7z+7m67/iJOKwtgFKZUe4mE9/2E1y4Vo7/Mg7Y
P1eIBoztLuJP5Oodawj1DcZFoTFcJgonjxmK+42ZPlM8Yw0D24sqx7JIp0FDZTe1XWXaktafFgmo
v2JOio8DrqHGONZAZIQPunaMTfn5K/fRG39vjQS0ZHNKmm4jvhr+QYrV95f+nxAuqA5eVQjF5eOR
hp7cZd/Edi1cYgH0ggpK1/TMDgjcxylDFGqJYbLVGLbif/Ms6y+bc/hjj1zKmihb/hM/6xtJr3NZ
5YGt4NUMZbhSylHAbpLXuSyh75N0RjWfG27kfOP3o1UdBQ62N7USfRcDoM5UjzswhGfbdxI/0z6D
a1V2NxLLym6ous/Ez1Cp5L3A/rMRx7FbFpmBqujh2FELIyGPsvGqbn9YM+Xt+2Eu3YurvXykwjnq
lUHiZIdfDRCs0J8Ex6tKQaT7bIsoXAVJIeYqThK1FjU+4RGMBTUhmC72Pde8cp0lja6RZG5r1Cyj
6nyTRG+A3d+d93B+fTWRrhTn3yOKp80GIS6uEk8glwCK+qqF16rnFT+pcMeEX9L2BX6XLg+dmr9k
CKRLnkhXMtaThjnBs+Wjlyl0ZKb0h2foYZaptNUs52I95z9O7pxR2w6lTQcyaidQPP8lWTcQSruU
ysohBwSNpDvBaX0G8Sp0+eZZSwER6AVns2GPqrK7/uwYigkgU3WJEPa0WENSpPG/EKRZV6QYqphQ
ZsjTuqXviOLW3W5PMRDQ35O+aTU3V4HqMEppCkfFDXzY/f+YBeEYpdsf3pLgYTTjzm7LOiBOPl41
MPLIjFsL+AjFem1vVome+eYJcEkLw0YQd2EltfgST44Z61UA+hEAF2qZdsi/IZLvBc6XqbwrLPNV
lOpO3mbi2T6I2q6T1xkamnGspr17THJtheWq0/TmPnAeeInywqBc1nPIsxcVBW6HqgNhuKtOSWKo
qlhlLx1TgyLXh0e4Tr1qnK1HJHhP4PIwuT3LxqBZoZEPIvuSy7T5zuLVLDRcS6rSi4smjKAk5uyD
3M51BcclGdb89GaHMGgrJaGS5fWJin1CG8yr024noVHFyXCEobFCbM/DyCdErGpYzGSN/Nu5eZMt
hmfIeyuwlmofstLgu+Wotalohr5UNfWv3+JV8p5+zj76IKfTEaGgZiuSLd3U466OZTmziC4bjKyT
kF/vHiBPGqQLGpDEYiMBxvhFd1F5MtvxjoxTS4exWWoRnFm8qMTRcylGz7FtIgurwdOK1f0DREW7
+Nlj7JMADjT9PW+urgjI/zr7lx4r04q0CjOQT7ndQOFVbICql2bZ6nnQFbGZx9bbG2ZW+rstaVCC
Ezpil6McU5YZHCEvKFxBU07gR07fmdFkqCjrrtFrL41ITCR0oN9m3Hc+Sy+ysSke3zPIINe/K+25
EeRIUINLZRbeSaFLuonrHoPZAbEDFOO6ZYwpcPNMIkhRiZFaLeW1Sjb+8AjGra8peLwgAVeWeQlO
ID2qZm2EjqBjvuKvrTiAoUpNbpvYd14gFsmdJcKhXE2uUPtmykhfxldIsnIRuLCX5GX67Wj027k8
oONgNEMXIvoxNeiM1bGzSaQ7qD9wZncUJlXnIwH96Y+cjIaedfhIQmz7JmjjwDlV3l53O1bgcANX
1VZCH3CothrgrLl38bq7ZDl8mf2ija5RfhP1G9RLZVc2DTNIKzoB1J7OLuHdluOWplRSmTDRkfze
yNAV5JpK983FmTcR5s8dh/fnB+aZwlVYnWSIUuwQQTf6i/lDbOqj+AqMtO+n7xS0FDII4IwHRQbQ
W31yN9gfK2yYTQXLyH5JcNRif5f6jTr9H2C5tyI7adfPJB9Jum3kdrDSr3gPYE1/HaTPPHvnwrmA
kvMZN3zhoqE+QJbTzBctupolE/22Tlf8YOYCld2bRAX7vlKXANvZ2D5n8vkVZeEVjZ/5DA4NBW8E
gTgExeB4G5vdHCpG8U23B1EIxubGfG66+C/fvspnYWDfr5UqBA22NTpg2EMNCsSKazYQGhzhWU6C
g0oFZ7cgC1NXxiafzHEERrd3D0nGDs6nFOXr+VO/9sT2LskVWG0wjl2RT0iv/Xg5nz+3KQYmzZLy
I5uiTJ0SIgQLuIOBmryfNQXriu2SE7mckdCYgbx5ZfOgofyXz2S1rjx5VOXraEpEg9pB4I18WeQ0
QlfdszYB3sEq5sTxs7zf3M5DQO8zJDnLY+IVvokeHKaq0m7bVBfCbymPD8LBZVeIpYwkB7RtyceO
vNnzFHuamDs9BZgyK6Mpg6QyG3L5DSv3t3XxJRHBbIqSLpORAOwnIutCq7XWAmtY2sAQtqoD5Bit
jiMB3TM6ZaBfcbaw3N2LeY+50ESXgHIqnscPa0ZjvREBIw24uwA/8Xd9VdH3Xi1UiaypXVQDZzbm
PJYNgoentisEJH/hQEonTpCInc26C9GjOvGxe+DeQ8d69YOFsMk78K8uGD7+fyoSX0NvLGw1um4M
kx76OFdbkMl2PLs52s9FvlTh4pp15bjtR3vNl30jPf1eBPT/WwEjVagyvzBNcIvrhdAN1J4zCGrv
NQn29OJMKRatKzOPzr+a4rvSI2YI5VY3xXNDARGTIsQjKBKM0Mp7aISV4fMFeOFMRwk6/iIrc4AJ
lpG4l2KV1CZpCYFSaHNNSGLiPM4jUJbbsjTakd/knTcLw5HzL2HH0Ld+d7WME03TCfN4eOoaT00Y
kWES151Y7jN7sW82rmI+mdLAIyG04mdnZvOpvLHisY8l5sODAylMx1a+hgNJXLiS1TMopwiqe4jO
vJPTYCz9mCsfYcDOhgDNYo0DbIfx0o3DXnjKTDIfVgO6mPWiXtZOEeer6nkTm22C7L8dd0eOQBKn
elvRJORLKol6cMTeZw1ga4sztfH8AgoK1yqfKE+6T25K6RgIKhsWiHrW+7lrTVmO4QJ0IWzVMkJE
gFfcM37xfl/JnkjL5umE3AcKhTbLg+TvhrWfWOmnEpyOU6YvRTjrCWouvQ5kD+ImSeCmotDZHrwI
gPClB3h9NdoGrc2RLZGLxAP/mE/IcGZtY7MrhhRLdPFSDnDm7kN/QPTsofqplVB6genRzukrGkcn
Yy3rBRx9rlLVwoMOJkNy3NwszbiK0XI2ekNmRMFowIxdVFbwJEGzZ8kKzIe+9j79ZglAZ78wBLKj
JyGsaxB8rigC0Yb9Rosj0qiKqh8aZV1cWHTG77hdQWQPjT3zNEJGPNUqAQwp8YTk3q8mzUE+f5cR
h4fvBduJPNIeN+cC6EPJ4xz083pFN1k9qv3mTaSCl422SaZRmbzdkhLivQYCzGiz4dNDEgONKTvW
hX6nDrJYrFTVLqFN5ufqvPHeznKwgm0IAAMYwarAsw2ug1mpMHdqtXSaVX5+l7fPfihXGrgr3FZ1
v8RX3ESM+vch5dyOu+U3++43ZBEtgRIIugfwh7rNjAsSNiu1tUIt/n3XaaAfwOmT8fppkYwI6VIZ
hDRoEnGvWFf3o0V7kCXTtEoqnGLS8kGanL5W2KPli3RNwfvTFxu5jB/wSQuKNMpsezz76SrrHlJo
pCrk9YNpuaW85H0514acWQYMmBVsUqlMtlP/Pyoz4xVqu4oFBTXg5NMjS9eRFO00uQTtk5tPpO04
CyklTKmYxzBsV8H4HqvEw8kt6DJ1+97AMBeBGQN9LLFmwijwB/nPCsHx846+rZsUW+PKmwgEluZk
2vKNZmc6QrrvxftpE/UjONs5HggAX4HdUfqneD/LIZVqFaiybfnfQWgA7YJncsgCMES73D4b888m
DoxTWrdartWWAiXNA0uTguBa+FSuxdvdIzHL6Wi/8Iej009crExI09y1U2Z4Ddnf+E4lyPier86b
07u2uyq7Z4s98mLlWrXh/ZBGe0u3MLD2VKvrz7MAi3bYoA6fpbVNJa1lKz1XZ74VGY8V5yLEXlD0
4VXFVExyDEToj9cf2sNsihswo50viNWf/U81fI2VLn4eg6fKYwzLdpEJrZoWdxsxi8IYp+NoFZCE
xl7uI9jGwp5WbhvL/MlbTGbhnqHOEdQTh2/1saqdaa/E/+iQU0jlSnn1CPJB3z8TKLbT+2h8BqRN
sIDyfylaHLCPOgeGlDXjWrDYVJ0Tjnku8i8F5J3bEzZxJsNcauFMqYfGbOri0g9G/X1F/8LW1rh/
Gd17xbaXT9DK7pRqwq+A9P1hz1GOw8uJtbycHolstG0tHYzNc5enTVw1bHL+lScUDIyOehLVEDwL
FpbPS3r1y6JDN7KLwVdrqEGzfA7Gmhcn/lpSLCtuPYwOQN6dQejZ27oxdsKNqraFojiUEugBCpLU
uhPkThfS+ROqABsrcE/u8Yv2VhrnWAr+n1p01L0gRdu1MQrMevKV4wACToE5Fk+lsxAtg9bKWxZW
Bv9wbVx9rS2ZLeS/lgL79xD3xTk/pcwMOUpUMxgxBWvJW4xBu6e3hYx3u13Mt9QHZ4ZYPpw2A1zB
DMaU0L4BKwAdN2B93ZCsQT53hNtxfs0jv3OgiNNVBFDxfj9nTe3QamnEwew4K++X/11JHrABrRdH
x+pyQvkCXNoA34B9utAHSC9O8RMg2Qy94AuIQIQ8gESdgSnSko01EsNOtjCAghr+qSwh0RZyxam1
MGpuRvfra1E3M16E464Nb6MSNlYFBRI15jjtL8ID1rFIjHBZxyNMBndaKPfRXNdZw7zvgeJtLLUH
65iqylOV+J3Zrg/dKPMGFmOMO8wcG7g+R87UaqNfnXqdFAISLvwI8FAcTeY4HgHO+nvD/lIQs7Sz
V7pgjVXTBDwCvTejVkJ1vf8UKhWmdnR7wp/Yt9sIQ/Gni2t+XH4Gg/iz5l0M1tJFNlm8VMLcHb6B
ypNuig20ITgG7pxTxwDLs8UxPFtK+4Zyms7PPgKuJ6916XnD2JFKxPehzpxxtKkNT4ASmb9YJ6la
IqIund9kcn7barq1kJHtRC6buyVLi8qXcJkBjntVuPX7/in3y+zN9jZZc8K2WbcKYXYiA67wVHcq
WO8hhBLtzlcVtaD+Y5mT1qLnTEyuWQIoHbZIq9axWAmhHTvBngsnbm6teUz1X0LPsQkDxQ1tpnuw
+iZ0T2NMDd7Qg71i9HVU9u72OPPs88Y7RD6GYFb9tECVLOi0/Z1iVEnIKL50wPXBcuZR+ZZjuqzz
bObrv2Ydv/UI9vwXXo8Ax2VdSlkOICZe5gGbZ4L+7tlSxPsUry9RDd1X1Zm0CkXG/qPrpflwNsP6
DWUbDE7Jn0Ga0mOPNzHAokq73+ddbpStzFm/9GRvjp1MjSts5m54KOnYlcLp/1KB3Rzp2vVAb0xE
RaBoRzs4zOAr4jlBSUcDiLPHaLWkcalzvpZYGCym41BY46aTKsGSV7XsgCPRC/Rc0fb+KMIc7FMn
qMNaYDUZjbFnCexFeFZ/gTqCpjxn/FXzWNPY6a4wJmT+Fd4tXtITCrSh1XcmaR4C2TBwmtKxviXS
n3JB6Afm/WHSO+vxnedQDvBKpRRrhWzPUJo15txDAsZ6xzrMO0mZBpdPn7Tx0mNN4NoG0xN+jdS6
Jl8lI+KL5RdkZZ9fL8F6wTKRSpbBa/UI7v3oR4BD/2AAejeOZs7VljsZ1xbK5NT2GLiEvPJ5O3Qt
X7MLApMb5YQdFzBRbWZCDlMjz2qul99Jp8EhQ4qrtmFlI3D7qRbdoaKtw9DR+pWXy2fV/3Oy0n0l
WdlehgGgJ1prIWKsaPAipMxYbHdgaDfbqK1mrYsgg9B06XF2ag6agCi70Txrnkh/qgA/3YuCOWAu
lD6eBMdXPnKCUum9urOXDWkhJLz67njRQmdXw7WNu9dlApb/spdR2nWIrl6D/p6ZwkcSrbw6hHkE
5bL+dVSnmuCpGNgbATKmeEKyg4RrbRcau9XuYlIy+Ln8sTAT4JnmotCtT2yarsrueVUbhDgzybMI
qK7QflkEpOuo5BScqYGkcGHURFGTXyG+6Zl+Ufg0gCy7rO+QI1oW2Zn7SSYHPpP63Xp0vgXVjjqz
AdvntPsTcUKg1RFXEISQBewpZM7FPx+T19xN2yaondSX/AyAJbcvC/GRxVfzy1F84QVdfMXZngNG
+tT6g0QfEJu/jQij2iNWCpuGykMcRgjYYFkbPjS8acASJOtaK8euqd1KEhGP83Tzd7n91KYJggFQ
qHhHnXo9kDo4QxMv40ZtxyBkGj8ONHMBUpfZUD8Iq44pwzEsfDtaA/NMRbUHp9DwFIG6F6su9QfO
rhTt3ggNfFk/CEETpmfb0iuTslzjwAizPA//33PHAmZAv9F+Od3fqmZIK6/DqEjkRbpVaf/s28JH
YmclsDzSQUC0G8yporpLnVsawTF+n8FsueSjV5ge2OPN2dKMdhtqVdk281oLCWnuYGhuhUvfxV00
5SL9wVP9f0vbTWLKVf3Xrlt02skdQMhsqegrU5iEYsIqvbhMaPt0gbQW98hntHjjulWguXwPbNkh
s0NNOJ8b8lVWiiVXwfTlyhEP4r5dlOSvRoz9hosbcUNwd7Et1HGgGbscXqEvgGIpINumJLYwd/rS
Tigw9AxBkqOtTTBpXaK72k2q2zsJ28o6Ekmz4zDAkcLq5jWEQzkKOPzM6L+Qa+OwrZ+EgM7n1/ML
F8M4SC4BK8PJN4lJiJa27a5KIeum8ToB4OvnIj2QwajbJkOsDP9Fc+3wwLd1MNQyz5S9A92YVap7
3AVshTLyOrz6GTrTCIsubnKrVCOm8JOaREzhKzhUr7m5mSX7IUddo+gOfkezBKxcpUdQRugDP97e
NSrNLUdFMVgJES4bxTp4gYgfLk4qfUGogdAJiu0gJlrr5Z/b0ey24lVdxSEnzsl++Lz7I8MlJIQf
pQ25p/BsRKSN2nKxVU10ecNlQzmvHpxrBiGrFKzFUqALyG1EYZxcSqT20TqzgEdXiXP1D+g1AZAb
Wp6+b1NGlPlcGfgxf329pAWKsBmLjTdIec6YngUMXsi7RNeWkNOfAqlkQvQNepgYAnH5Ks50IGWe
CAiuCoPRZT9uPuY4pRtr9SnAEtlYJ3rE5pC6H2JLKL1OvTCWrQsKfm4Ezz8snj8x7Czn6lK3eE9N
Oa1ASR/A7+q328G4oKE/UbMMeHXIv5qdk2l4s2HnSBI0kM0319C4rlZVdUsAtRPoODF1HohaWeCM
uoQ2Cf+NuC8PIgx83MoNxiQgntymUeDIF2AfXn49iZMQPkMHghfx7iGky0d0rkD+WZv2aN/fBvFM
loMX2K/ijxWIAeWo9bPoKe1wG2YkE7/QsjB/BWLIlNxn+VriRn1FcFUnnjXlZGHK3qlXY34Ima93
3koDw9Ih3mIGhrM+Rq8mpAGruHnSOYxHWtNMLLhALV0ClRWl1EZKRKzzMTBQB9gMP8haabbCILtl
gVsItZBVOrVvX32AIHLP24eAdLy/5Fpl22HBFHLXSZD/Vi2X+AAgQLSFZtDv0BeuWpx6z0KK9wPU
JWpmI62ymt6D2CL6vlpODtw2BJ/Q/BTMssuDJ7RS1K//IpuO9DiOCxo3F2ew8xmt3fK3WEdp1JFH
v24IrWe0kZRxz1+xRWGhbx/486tz3pFofo9NK3uIWCIEFM5cGJq0zZZ3vE97qIFW8pY/qPtCB0iv
fiINSaxHK/kV7XcoyrOxETPrMqnClXdNJSe0MTAfl4kyx6pO/mmnFS/ej4+Or5a14LK/y2c/2m3y
rr+3eRL9A3lG2BEPewj8DlQUBKGOAxfduNLjx/5hD+/0jFKPbDMVCCNiJOReGG2TtSQ+ZspQIKIf
ylSOcXFA6RDLlCTr/72qsWS2mzl8EEZlGFVfRmyzdMZp4vs/Aynt5ujtxK3bKqIxYvcmHt06ieeT
lgDFgw6mdF6QU0NE7DZbWYRgt+JoK6PrgrxgTyrpJDARJi3cC+s1erApKPsoK3lm44qv8ZtxvXMD
cFskKLbZIlR/ZX1dGXNQpnTSm5ZI5mwwIPt7EwxgUY6XaEG+umqV8wSeAg4nfKHLsFQMsqRVqv0R
58oRWAvQbnjVa/WVuFiDDKG0jt4HeVpgA/MZ9DS5Yyxyw22Gv31TuIgLdvfGLaqC9Ua73OmZMMJ4
+NYIs4JoMNiNVsDkBRIyAUwJGh+VvHe4A2cV1hebI2Z0mZ2i/cyc2OdYfiKUQyF+sQEhkc40AZNt
zx5GwSdCo60NIT4RZIaifVeGI+PCnsklVvWLdYC8gz8H52Pv5OOck2I7Bkh1JAsVCxDtbG8IpFxc
KvPMtYEGQl0cqJ1OFQZsKAMR4JScePlk9sxhMfryyqTWO3KhX6dKwl+3hBvEMn87kpbP1UvrVB8K
PfddAUcVVnahN/HyLijzYit8d9I/6NVZvNQWOc7KirzYrpbRhXZf3JqaT4JSWJeyjbUiMqWsa3BI
mETfzUpTbk5zwavtysrqYIiihI/op2PRbho4nRH1DyePJKV8llPdYExxGfPIDoZ97+KWsm8aGE33
u7L2sfqc+WHiIy+Tt8zHcsQ9ugFlGhHKZ1LyiPPI+SRCeC06yKi8z/Z7FFFeGUxXY+UikR3WgbsJ
0xWNPANSW07YJxxGvWaNzGdnhl/cIOkZxRdYnNbPyf7UJzc3bXzACGtZ61AennPunBX3CJYphoAa
Dh0wkHgCXwqpbUhecIitgWgVlLqrU/dmftcTO+Hjj8Hb6UFxM8XhDBv6uYMDOz8LxZGLsJUVWreu
gDPwqOTxbyI7qZOT9TyacoVMI6g71Xrvb6OgKlpuv9I0urpCF+9zjW394vUoNXUjkx0iFtx0aBZe
k4OmOO7aOdWQRBNJfSv/FxeYu9ndjTMX9NCbAF/QlW4EEB3a76M7pCs9cr0r+IN37Bo5kkGg4Th0
khpZGqpn8cXi7KcQJFzNiOQCMhlKq/o5PZ/WLrbBv2B5Y9IVxUYUTG6k7cMhKPZvP2EecmU/81SA
NSsgmESMR6jRECYo2VW9hfd94qbaNehJivkslFbfWmhP8gxbdvTgxWqH6NAzmKmVs/MLViaMQ1xA
A8zm69XdZyzSBpYy0ktx0hIcnkMQF8Mcoc+ZwgN8c8640EpkgEyHDcOXZREkt/x9klk8PfsZ6Xxx
JuUZB8bA5RBZ+FF7T33HqR6fuMCPs2PQde0vQ0mFbIx8lbtpnRfnQ4QwB9nLyH4RY+LU/XNl7zNS
f6bwIleejsrJYsCxqtCsdj4he88+WrbiWexHcb8TgKhCr7l7SlMmzOzIF/LtL/a0wns4n8PxXfeE
m96UpREI2hvvBPl89EfuUdYaT0EUJp4g6VCJfE7ZPRrq0+O5vdvelRtKctDPB0tBdPFEtH1Dd0/6
WpJirIIYIB4PcwPfBtiQzt/CGwZ5Hnehkq+ze/40yTLOX4IO+5HO6o4E6tbuz2zRiJHz4gIILhdB
1C9HEDVGmKcrCG65aSv0Mb9aePOB9Ms/9AY9OTknYpeJiAl5qgTTcdHL97/PL/8Ld1b10NKWVSlK
pCmsSddmzAp4N9IK+YxEAgdCkLGrcd6u4PIUULwndCG58AyjyPmSY2KPoTqnYVa3GPkhwClpyFZQ
lGGehybt4H9Zg2x4IOAJayay6DkAQvcWThECoeA4eyhTlUAAeCUisS1xBY6xMjslb6zqo+uwOcE+
KeiCU+hE38qO9PQY7+91e5wv/1Z1x9xzCYQS9MtywNwyRadH/kKG4QrrtD6T0gKRNDSOnP7TOL2N
wyXwv13hJ46l8wGBHNKRkkT9jQPuvL2dE7RodKNmw1XGjHkElXz6vc8YlQJthB1vYSGdkVt7AwqB
1zEyYlHSFWN2hfP2379hfP3QCzppEjRY4wxYNGGhm3FS3yaQR23j3/bdYmTgF3VwGR8AOZL641EG
UYnCYr6ESGsf0f2PraXGW6Cl2lxKXcwr1GXV/E3x1oFY+TE3VFEjuOOKibLzF8uaFmk6It7BXSQe
RWlMYEJADG+RaCxYFYUekUlZ6jBKduD+EsNhPAvsIbGETgP/1dE0IEv2JDoLnhWwbwfePAqT1yke
i9cBNxDGT8PkkqahStJw9VhkBgqlKhIcIM4b1b1n2kHjxfcLMxQMot0tAHIZKfF9CCBg9CjPw74z
hEMK/wjv8ilACJBLqK7FPxYg7iL/K9B0HTSMjFIeQ/CJfn2PbH532xgr59fRrNCBUPxkxyI+CPT0
xiAC5ghbU3VHUWr0QrYwxxYz2WG1hnhlWKc1NhWoan0r6ZCf9zDiBnRUg57Sggsh0xJUgtLNjy3S
iZIOouLIm/+n7Ft3FVK6S72FkADGc6ETaVHI98Bolf+OQIsBYtLUZZrkLbxTch9zpIfOomaS6zdH
92di3QZpoNipCJXY4Nl6R7vVoLCDa/ESZwzGfoVPodxNLxx7Xx4cjJ5rW2V9+cXzztIliMSk83n0
GqJ2YeWfNhX6Szmiqm/E/zsjP3HJPdVPD9MLE4pZgcq1VVcECCzuXU8lDC/+fzMatW1i1RoYFYwn
v7y0PvDtF+D096eLrY8EdUnXQviMWr6tUI8Kg66WsGRJgu8b7weykqYtsSNQ4JeZ/+DMAs9MaRL4
0JVNGQ5vIygwzvhGvmVJIsAAgEkSHdAX+ZV1NWC4BXxt22xTN7t1sH/dZLi7kczRAjanWYHm5pkJ
bAcEACcJgrQDEyfERYocFLXMcLd+JN1ZWjxO/AOnAr3w3UXiu1P0sWgApWHClCariqGUe2xecjLA
J91HLcDtXT/pr+44HDKiYiZHROSfFMGooiqfImpf5USVMCc48x76TZCzfzrK0U15VEc25If3Rq58
eZ5L/ZeczUIfNy9uDk+zoEHI/wrio46/sJGMpzzO185THPfXILBMBa59yWcY2yWxhCr1tlJdTYSY
92n+BBkqGSsN+P+RgtiCes3uzzVwvffAbjSDDHPq2oMUGFHZSK7YhZRN1z3KRWTvlPETEQq+h8TS
xMnVFHpmA4usaXoKs56jtnFTJABIZwyNjIq1BmzNI38RuajUlQfxln2ElmGW6oBDpnS30QTU7sAd
/HqfWCfsMhJK3cz2Ux/8JZJv7B7oLolHb9mpx0kmMxK7szZf042Itw3PDZoJfqEO/Hv3zD/lmAnm
7wHIJ/LpNYR+4oqlrhmZmGtNfJkAYVVyY6BY0XME2xHf5rM+8jVD78G50wrW91zZ5quVCPbtiqG/
BSiJlPZJoM1ZlanKzivR76Xt9hu+LrA6N/6b17bltkof15KCqMhhCedjeg5gEycxQkNMqSDQnNvc
Seg/uzs619xpgn9IWi6jsbmdzcumrnJl8tqbJ52ZyB7nR8JVre9V/Pc2zb4pDmWUBQpoSQBo7Y9N
ceiopXzjo78qbNAJsdfl6FEy1smsAU0LHARTSuKkd4V3gVBDP28s4ir6491MO7Tbw/shjzuZ5C2r
GaQqXLXSPjUvO5DCdgaTzMzbzZIhHy6V8554sWaDvhsYGPVrbP9GkjeK8IPGUWLE5kpnmrXBGdID
RoRjHZ0BNWwM+Jc3oqgMK3+42608mvuG54M++2G/oSDXBfuG7MuBiEfX0iSmayO9EpkCej6ik+TX
/I4VLEUbW/xSeyBUDLc9xtycbJNCryVZ5+hvEJQ4TIyELyy7AKkpy1C+HX4WDkx11xK05vy2tGHC
vjOtAtG/ITdFE9ft27dCi4ZmBE4MorJeAvT9+jOthaVnhOLC4m0REHP0ZN7f97hii7pDwvabT7gf
SkZ/f4WhirTuX13fKWgbC0Nxu0BDMX4Z2G3542UpGvMMRE6Ga9ZusRWrZ0A7OrHZ0sE0680PPPY5
pA+dBt0XEO80BuLkkD1lgermFohvO/vXBj1YBl4ZZpwztWAiWmC5VU/gBCfNFLYcm1hj0rJcuEK/
nvGhmEwoOsSIh+NMxeDVS/F6IZ051n3XcmAGZA2J1zD19RBVL26qAm3Zm5F8wDPwaKkVke7OVxrH
I3MycfJNg2Hkbuo76H7HTwrib+JktmO2pawyXT5oGEndOSX6G+ACyzUD7gTkiLc7urR1qV3IF4R0
7DqKBPxmdLxhAWoZtDX2YXzDyKw4yzUJagnmIjVPtUykCMjn104Jhi1Zz3k6rHxfZIZ2YwHSk9E4
4T6OTXJdAfTpkQBnqA/ZMlzy3YqY32+cLV2NuTC84euYSw42p/tP7HNlHByZ3ko6oSiieoS8Mexe
YHqaTlrp8uomuhdIgEXkLa2qzcerxCdJJUwXYElJbyC/GEBnWNL85wJezaR/5SKk/ohuZFWVYytt
nwRnmAob9t7lBo7DWQRppElf2lnPR+G+Lat9TSsjgkX6x/NTmUS9ScqgNH0FZVJXHwuExbB9BHKh
1RwPqUqaqFiKfcoXaDPnybFublbrbvuHI2qPqRDBet9DX/i0i9xgiZQJymgzcIIEBItQKhH049lh
wenjEVQG7LE/1T7IWTui9rwM1CDuo6NNGhk/pPDEzHr32uicOFwjv92aw/UeFZODrBZauz0KAakD
GdzTAzJkLgcaif0m6Qi8ifDt0Kn0+eJNDjvKqppDUtZtFyksa9E/Xt0TtKDRdWlzrKl8YZo0+dWb
GDWCTBsPWitlk1WVTWp9Z8UnAiZnlA7ZdpJVe7KAImqhi2jeBlkdEQtk3EE/xdBmiR2Aa+lnS+Zw
c39sxBoNQ+pV/D/LkLaf2UOJkEv+XZZtvF/f1UGOiLFs/TDuvAZ2e5j/lA5em1wZbwqovf4aFkrD
PeAwrQF7CnhtHoeVsMqy1s3lyK2SyKlD/sYZmC/kGK5V9khvzmm63cmbZWL0MBKJMvyPiqhLAlyH
RBRn2gC1j6gxbslZT0QylpLcEYB2sN66Bc2cmjZ3EASPpd3SlxSHANDaqZ92BUJM4DGsyi9eJgJN
tjq218ykq2DdSEgufzhCuY2+LxEQZmeuXahRERSNLJxUpnoBltArypUs35piUWfr7I+1Td1oaR4W
GD/GUb51J0194a4WtCE2TcsG7fkib7jPAXa6dqzlDxzSp56KLavPhvbU1WisK47myRd9cE87CF+C
M+C+BZFoi+ehPiVP6skTTnIc5yFVdLabnAf5KMA0k7Z1LwNdM/dWXYIQMlF7L/KXSgNsVFwSWXAQ
NgQXnPH3WPUfyocrCbANbWGPEW+ROxb6OFxMUiao6mg6/ywNbReMHKDWxOvhlbeolwRXWuJPq9Hw
Z0n6z6m0vYaZJgIkLCRZQd11S0TMxoDh38t/doAAcar8waaGyNBh3QNs/q+/Cl1YZEnIpy+wNxwl
IMd7e92AN/0wAaq+lmhD+H38IubIdoaepHlot5OTu1AnBy2N+377gDvQqPOTeFEKgCW0Tzi1FUYP
ZpSeRm98N/4ghCU6cJgzBASeXlgt/jBGkj3MJtb6vIb5Taq14vJyrqBJ1xngi4Ek+ev8XeG0Ro3p
nanQQx/7QdncR+hkgnKfSgArUS2m5ul8IL9qshcjKfTISaFhQOg4omxve7zilKaCCoG2C1Nb6VK8
f0rgHkIPjkFnJ6hYhOElrmGwNpu4WuR42rqqBVeQqngVwKwEGxRMSXDo2Cx5CZanP0AZrZE62BdL
wLynbEc/ImA6LbgEM9ce1fuaLC3bYGsEWdpzU6Pvt0DIITSOL5JILxt1DS2nYVsBNO69lGMEq7tr
btKGppzGWZ5lUmBxb9p2wSPYl4TRRSFrY4NN4kWoQJLm/BeaLkIeilBXfN20Ab89RydZ1NGzzChY
GYRGZXqmVHvS4PqB9FPXs/A8/xy2Elb3fBb27OJSAKRLDH0UOVabwlIr0I3iiVSCm1Adcoe5fIZe
ej9j9hzzu5zbtqOC4UCpWw2PYTh08aFYHeMBH3OZkX7NxRtmQXcVrmlmpiURe5nWM3MnSuF70miR
9e3KXBSy8PYr/ceSZG2/HnTs3nJmu9q8HjRZfJJli1djsSzPSWO8/82+JOx8AEYvwp3gMhosOMzx
r1917CMhMhz5NaLQJSROnDn4l6bIGFOuelw/UHSAJIEBzjvxzF4kJGf2sySHspkeu9hFH7XaV56x
zlejuJnGLvG+Rng+sApFSrk4c8Ga0DryFH78oGQ1GFoCQptaDioytwoMesmHSxxswo0YRmAD7+by
qLNzNTQ2Z/0mqb86DRDDpPbj2yT0AaekrCQ5MFUOorrJFgO8shRIzLEfHdlaAsFZ7C79kZBvjr/o
yU/1DqO6OaJ21PPqx3mA7I7ifDj+edpLTfJzuy7LtK2d0RfKM7SzFYiKGZ5JjVhj68FzsIkYiKYV
Sn4/d5PBZn4/JaylkWWX6c+hEblxsKYltfC6/wcTLRxP9BaoYGPjR9vxmq5avy+2O2p+B7mcGrh4
lPn9ZiV5IYCqu59knNW13jNNQDcWmuivWuOFm+46X9hYTYI4PUNIC1pQYLery4TF3ZWCOwlpVcbe
gN1eCUpRWLYV5fggv11Tmq/vnvy8isVN2HPQ8248QrFszXhD1NwpaRT7z8pFXMt81VjlZ7TsHUU8
pjgfq90PcdeV1E+Ifp1zgQ2tuCfgtwg3X9XwGzWqHNPvm99ST2PCs4xgUVWfvSTj40GzlnK+M5US
IRiOxfgIv212qm/ahzHYpLTcGmPnCuuoh6mRHTiTNNdnR67511+f/grv8vvwhaBLlTHJad+el2gZ
j1IdJvrgAylp6ANLaSvXAyjEJNEW6r8tKaDRoTxytbyksgELEo3yLbxmAPmmuVEZ4nl11BCd0qZC
B/iBsJ+YoGB1QbAgn4RDkBAaT1ruVRi+WC533vdloOqIa2V2+v3C3w2VItEak4YsdeP1rREd9iM7
AYuBRFO4z/WjZWeLK1WIzKOjWpFltRZrxAl062ZioESbqm3hCrfvom1mqAnumUFLYeo5S+jP910e
tru7h1UPPI186SLmF9J8eq6FpB6D8hj7OdgBc+uMIOrmSY3SyXiLht35MZlyCiMBqkpb60jyH+ne
Vi7jMtJxZJqtZp97mQGtpaJBINZOcSY9Lar60ziG5MEEezF9hvGQenganvYdzLJqb5gVUCnnOnsM
Q8+F5n7VABAGCWePRnJlCgVpD82igNMBVId9eBOFgQgZlXvVbblcq4I1hIUoAfqOxEKivZu1XYaZ
lNRao/i5NMEDUuP9woGUbcW+npr1Vjz0+UBahlkRk24/UkCJSSmBDUQ2IYsw64317miwWXAgbVU9
biBsdLmGuzjPCU1OBf8lAy5RZmc6YJaX4Ho3rnYXScLQwULfVUS3Jfwm2VmaMuiMb8Bege288n8S
98Fc0x91qw8+ezM0lwrFN0/KIomy9oV8LDhs2yVwAyZ/QZzwrtBjD0xtj2/VkeaaZ8HOAY+1K6jq
/nzfCBqV0LJGArdQi55t8tSeC6kV3qJCufV8soJFJ+8B2tsERaldAovutFdm8/AYTE7mj0u1r6TS
pXLztUSu5UVKp+gWV2IjA8T6WuUZzrF69PDcF2eJKFwFLQ/hJQElUq099MU1MhQ++EOnnm7STl0a
5VLa1I8w6cPfn8Yqgs5qDhCSguOfiRatLVRqb1EJB6SDgEC6/C1cNz4M+Is3x9XdKK2vwsQy3olk
p/dFMVnTuIl3fCLXZgN2nmrU5H7g6/IeK282z371MrVwtfq0EX/7S+PIXaIdjZtxz1WzkS2K2Zs9
IO0opsafaLjVR36Ij144hUfVZZXArQp6qNzLieGGGQJ/U9zkb3Tnq2l2+MXdAfl7RE7mc2X8YNAf
P3u9U3vBqDbyhcbr0PmvBwviFjFSmf4WkcBu+yEvM5Vm7LLNoY//aANcQQvKUxJ55ku48sRQN6RA
IVrw/oWxwxkhOZYovuCoEVw32W886+1snz0wqU4z8ag0Txc1r7p65tm5q8Q1NAypApSiYUz/FTc9
ljdHeqYWznlxHgYE5QgSrV9hfFvZ7JAaJ5hPYon2z7sxmb/811rBWRAVWXFB/5G5kgdGA8oJyp83
nbc3ClJyGhQBj8t77PKwv8iL8Y0cErIJQxvXNs1W3O2kqlI9AxKzbePBLvkxxfDrKKPG9XmIqWi5
a48L4XZjB4mSoMoNXHAYhL0xdUhpiIpG6left0vTrC4SLDVbMvvPBYFJNA3P37ZwdVoPxuGsEE8M
KrqwTCE+B5oYziGEQY0zQomuEZMHUqSgrUNejHmlKt1c9pl0rG9BuXK8YlS7thWTFcA/bZpDnuR4
HN3XXa9wuCiEbkaHugZUeVUcknyjcWjVn1CQJc0rDbAJNkDRgAQylh6EhTyssTsyFcDng5KrDM/K
lXL83rSa35VF+ITjK5xz5jI6bX0DQeYdwvLzSezwoTSx8nftrisUPfy3yeQaREJ+ybniQ5tiX+Nf
uAhbqlHPsNPogvxA7Nz9Z/HLn13esRjVFjTzC9boKSAVxv1AwI++M//+OXW/LZtQoUEAUDYVcGtk
p+rSPb12gAxkpudyhjRf7eY4ho+SPgd3P/sPipFCkJmOi1VJKM/D4LWSqWdSabo0eY32hp9tbFEJ
mmCmkA4yY1bJd8hf08y45M5TCCmYyRdD14eqQX5xsb6a+VlauVaZlCOy+2fIbmXCGWJQGfIrDYz5
v1xlz99JAgJgOum3CaRSEVTyPdnVlXk8C1pevuggGEwHOM7MXX0BwgURDH49gHUKNZHCQl8B7AVe
h1MBctNym55kLvnp9QHF0SpdSOA0ct+xO/VOWdnXyyIGM7iuFR2+J9pmZV8a1QdGnz10ijUCWo+b
I/5oe8ANR/yx6CwEwGFJaYFXqy1qCfOeasa6ps4orU+RSSPUix3aLPzLuPObugcy/K/ZjW2XIwaw
c8visr1raXfDWGSXqyppUk9TqKCxHerk91sjShlQTeLFqVuZfuEDrLmLKP+oGyjs9kgL7C5c/Bbk
vUV39aqaVO4K1ywDaAsZ0ftfAsgYIR9ywEbpEKCl+MgvM4WZwRz6HssCLtMoaEt0ppns6P/KAXBq
RDl6FQpF8Or3lQwLQcl3NSqQ6fbmS0arDwRx2gx85j5vNLH4rqom4lFT0d/b2VrjMT3kOMF0CJa9
dNeEYD7BheNdnEhzJkXrxkst5jJmcKi/R0pBgjOnTECRrMV/2MeIdVB31p9kXVkrwUfI3oDp+22k
UMK3Iut9nKunuAoD1XQQmCFTat++xafEkj4JkjfFYQtGWjncFzLqOPJ75Y0Y2Oflcq1Iar+NoDBB
xPCERNNd+k7x7yjLVjQR3KK4dre2PeGLJVBh4ytmvQ/u0TesoBHTb9xHz/hVFZTQ6rDLLMdz4Jtm
OovratzSPRbwzIrejID8tCOcq2OMF01FXo78cCIyG1X9/zsO4gEH4V6lQkbIMhFwQ6fgaAKUzyId
EkriMphXpaa1Abq/tAkNoj9vpgJ9LIl96vssP2jQmHdmEIxMTcr55d6ygZmX2WMgk7qmak37Ba0s
4LRTRyCxCKbuLGheVaGr0cs0AgY43g3zkRr8wXU+0tT/SriDXVsPN/94vS7+vwM6x2x1EvS1yFU9
kRR3JC3dY3OVPFLtESvE7PTaTEhAW9FgmD2UmQzeHYaMComVEsrJzLw5+h0jOt3LPxvvANKSOVck
muq+T/O+zD4LJXOYbClRrn99otXDmC5eIcGv61tOZr15v8hmVcM4T5oy7YCSinffNs4PILojTGkL
s4+zoVzKn5ExjWCdkFGY7zbytYKQWdYxuyEQm73ZNFn86x49v4xJa2fbmDCLOu9Xlw2Htda+QLEs
YBU6H3b3ENmATuJ9NrEZiZrq6B13ViWThAfM4FbTc/wIHcO0pJ8nPTx0um9pUE8WP2RWASGfmEpH
jHsp6vEScxIiOfhcGcLGga3uK3R5xJiQfWcxldKh4qHfV1xfFVnoD122VhE3YaAD9UcrafnXj8+O
BFYBlMiGIpQj5KS2y4xNZXCWDCpHLLsIMVrAWhoSPLYSRvjUqkFLH+C55OfNt1/jn+JHkGGxWfSM
t3wzySjIlnGycoCvRTeNfqwEiw9lqYBHyNN3XyXMwEfbV3dmxzwYSEW7q6nOjLjeDI0lz/rrye9G
+eFO9/ZndpdZz+FuA1ZNYUyvV8w7xDzrYcgTydN9xRuazCTZyT1KDoEJ5PdNsXnje33MR7Bq/jJ0
uokQ2Fa1t/oVKCC4QLMIM1WA9UyIBLF38qEqq3hJYvzicz4YaRnOVFZXgjsfY7AkcUIMLVWuzgRz
ELZYqqinQaR3pFmREyzQthq3TkDU1RWAAmuihlgcDafMQXRNv6FE343aX4SJqqlgpymgF6LXHx4l
AbTcp7IyK9fzST/0anlNy39RxrqTD2nVvh+IefK4/P6SxQfh1+K+fnw2SwctRcaVvyZE9DEkbYU1
X8qQHIi53h1eak2hUV2X9BJtXjboydqeF4BssiI2u/RT3fV7JP4NI9L1KPQRzX+Qbdr7tMNn8wwl
vF0+FqRLSPmhauHhXl4DZBWlUrNFRWQGXoB3v6IKR1phlfUYbloJTD3ynwxC/kedDwFIcjrZFEtv
V/vEVqvB52niGGHFtpHDSqlbcrpLbrQy3/upDQSPmhKyRs5avWLKEOV8saWUElt1pD9LIdf1E7Ad
5FT8Jak7l4ub+J+CXwyivWuEMRocLpSS1ItWLD/RnM0Uk1rUQuuuaodD6tViw1eipjTfvPLFGPY/
OpBS46fqFkW9opA24fvYyg7DgcQfRIJChUKflanNNe3IiTtllEwdBosFBASZRd4ihtdqyeBm2swk
UwAMkMZxdczJ1yKZt5P8opsmZ3QEhMKaxc/0OqH24Prn5DkiUqFDvgzRO3Yfg8csCFjfGpuxz9Gs
+I0BiPdn7SOelnUqrBJFucb47d3lMg8r3f/55QQrLjv2DM/um8Yep579xy7HBK5TwxPLYG0w+tSl
sLrRy3qyik/co0CXUkH4hLM/nFWae9MjavAHS2UYX8ZxlACnsDimLsF2jdPDtfKMGyM1qxyQSMCJ
BY5g6xTPuDpuDce+JeYImpEQoWmtsws6/KXXYqJ1qrcBVataF43HW+aGBufsvX1ztvKFFznRnoAs
XY+qA1EPdYMMBG89pdr8V2xccBMbH46uVJXQ9GeLMU563taRvnVa33ViAYSgulpjNHri3RKJVqEd
4+lWCXje3AAIbDHCNbpqTSkwq7P9s1QfIQLlmla/nzt3oJfJ6ZT6n9xtkOSxe4m3nBS13MazmVDS
mAa6wN5KN/zZfWh2nOQ1J68jhXpsKdr4ARC6yVex6+1xNJMrYniohMDi85yVId/fTXgu3Xb1HBwy
jDnCB/RHPwth5u7Zp0d4sv2bF0VQIysQM6Rjtokwy3xPeC/cfpZuGAW0/eJZirLSyz1wFiVSEFN6
tVNe+vYw9A5fIAIgO4aphkryrz1jmgbjx1Wbb44SEhu3MMOU8J3gOLm65zDTG0QUXbMlTOwitq8x
eIGmboeBA/7ThkBdmRyan2kajXa8+9wlOGkoEv6s8DWsuqfGxybH4FXba7sQnGZLLY0T+ERpBghX
77EL4ThsIwV7SOqbZWZk5zyDeg8KmUAuJiXMpOpGDXnENpttaEIGM9yXRQf3q2sxvn1GNp4iTNHl
L/o7qCXIgau9BYlGNS3oWE4W9SAzoZXg8ia3rs0GaSzGDAaMFJ/Y5fp7DUnrkranxUzWdAN6bFC5
Q9910vzdhSmGrNqegUaXT0Z8v8Y5QKZ+YThGc5i1zpVGh42cKTp63OjYLiNb8dWfi47ygsB4gdul
0oG0VkUAIYHTV41qq9yed2MvhbR1GLpAZ0zsoMBXXh1EQwI3bDmio1G8Hc09qIlz0T8Gjr4/yebG
+EEYaSa/dHJ94mBmDy4bUXd3eJ8xac+czek7HibzWChzPTPOvjr/BExgrd3uo/7WC07V2ogU4oIO
z1a3UPCOJb2SAsdwCQEeIPG43owN/LLXw4jkYbXX0SkL2tQbVm4j5pRytAzAhhlfP21ruU17LlUM
2PGGmVLiaAPn9FjyRRjlVokKAFodgjyCQrRhprBUYjt05GedG2sTmCaZnQXr3nCIlbq6kMdpdiny
58xujhyk1bjqP6W2B2J3U0sOgbPpuar/hx/td07wQ7aUsos3KPoojGKIMTM2hJUFRhIeDGPXWdUM
OjbXKlON76jh6Q6jUkCLxzzdgj5QjoHvbiwUkydA+BIjzvlvDxcUUOboTP2d8s6/zeMsoAjKJVKx
LM1lyw9NLuHT6QpSHrXjwi9GBBqffPPbxxCeB3OXxepULM8lbOfX7VWve/Bl37Y9UBCh5BA6Xa90
aIk0L1BypLOBcNSUcBl2IbGmGGPAm549oSKUubtjbUBYSyZt56/izD+eat1OlEb4+xUvfihZp6as
81PU6uzSFNcFD1B6oqwGfbDuTbVPqCRWZao5GsbmipTqD8eOcQ7APeT6IxaiJpc+XARbplBa6FAH
d9S/2e8RUwLhX6rL573mUIh3vyCXeX48mb6pxPTJkWPUMCAke+CPfk9odiUTyuAB15+3duHLX/sz
4CsgKPSzpmfSqSvfIwCDZKPueZAk3Bm8SOWJUuxMapDSQVgcLugLg/GkKTNZhgnAs5PHQ4RiE0vt
43qzbXVXZvbzwYboHKS7afzbJiAhwW8Xvf2ER7mPMv+QvTu90C2vBuwr2QJokLDouiCnlMn5aEzj
G1pQmptgzgg6SvCzo2Hjh7ExaPHDJk2lEldHn46fIw3IZaNIhd8evZ5Ja1d9cCd40an32zn7NYAS
Ur898BqZFODnSbk0puBFP7l+fmoZEE8U1XwC6yNsgkeRYR6WUC8rKyd061gbPEnjQGET+MMZ7GSX
1k4TGLI/cLIxZu9Ji2OYYTtsuqfFskTCmnY6w3Rb+FWK2Abc/qsprQd6SUWx5AYV0WjlxzNPtBsn
UloIqXnolpGmue/HlWO73mYEoozWGILuAaiJ21u7h2odUrJE+MsdhCL104f0VkPXfBbFN7XHWE+K
F3eJWDs06nD1T9vgf/pg6Mretf36XW4owArG057KF8yq5Bq2kuA/+GIbIo1EgR2bmO83a9Jy7hVz
WhXBxNYfgXHhd7p1rj36tFyELV1se55YyEq383EvFTgUCYaxvdb8/Il8RH2LXrWzOsKR7X6biMUy
Z95148/2V5p3nMSDzKZa9ReoZ7xUVTYb6SiRBGl4Y5oUrUtYmVfXHtZojTnZsXFO8Elpt2u2hH6I
IQclM+j5mmmijUHQDjWT3mJNlp9caHSGxpKGs3sD1+MIgRtg90dR/5bp2aaoEhNutP6uYjRGXBDP
A8HRfD9psRIQ/FG2319l6RqqEZCPnYukDU3fPVlfbNEUoJJlC9ITBOZDP7bSWNdGCTr+OCNZaPeC
rJGfjkeUa9eD985qU5Pd8alJ9jLKq1bTrUbPArOKY47B0yuUjT8/6Jevjlfyy4N5WmeuzFcGCllI
dF46B5cPY1Q7Gggh1LKNU9BJyNzxHHvC3E8dyo8yocfPUkdxP0ROsHCwqJwQxkChS5cYzaPE4snV
dM4opiWV8t0cT72CuI9A8rJpSV2P5sga+zjdbMztX1i0jAGx0lf6eUZ7mrYAaPmLy0hBMHo7uML9
ozZiYbYZZDBGuWphVolMLpiSGmId/57o7vfMsuXqlqYINKG2+lefpUfX8YmtfFl6AG2+PWs6cY9H
EWWhy2SMGzWqj9Q9+OUqcepr7OZqLstiIZgPyKA+1ruSff6H7MzLZsVvA2x4B+aXH42aioIuqcm9
a8eF6SCmwgneNVBjAAbju/oCx5+umhX9xO+fhAITjnJYnmxgwfoDb7QCXLyfEnDFlkCOxEZtJ+2u
AK3p++CuT+YZRidiQNWEfwdeyRMie4FaaVr/I1zeP31+S4UyZrOvnB4WjXjCxweD1hKx5pt/pSG2
KKVuC4z/DQDBejkEDkdnB9nVyjhVUHV1fRUiyEOWfihkKW+u6gYKmC1Pm93BKS7rlDqpEPD1F2mP
K0Ln6BDpesBWomveqKrzBcvU8e0nT7tPN4TyqMRfQZ+LyzcyHx0VvtoqYLYF4bMtNn0Lt7g+bkGw
C3zSAcbxL21xbX/w9QOFm/ee8IJ/i/XNKrPcFMuxRyfDnMAtIbjj7pG45Op/WuCyBQ6dE8FIm4xL
D5NV7QjLDjw7nWakR5xPQTOLxbzdP5fP+T2GcLVyd5CeHZ6YF5BjojMUpEIiK9VqPyccJuHOsbnW
Lgrb2FlvrO1UcTuGdc5b9CO9aBfWaOJKbqcMD8uzLYfGXwYbFOlp2uv9ReFX14dIDkh+gKZOu+j1
jXSO+ulCJvyX8DCahrlpLsqSXFkWuhrCRARCo+pSKmu9ifqvgIfHvRSoA6BFbWfLC3kpLeOqGKSj
WCIeXVQY/WbaJAV43p+U/wR79j5sySKZfApGWsX1u9fUUa5ShIYU4nSuL05Etd8QWi8ziKDPqcfE
cHVRvWF7j6sAXdvi+3BU2GLE5mSRjLWsX5wGSnmPha7HKzIZrRRrIaMP1fqwsM3wx4tV9nba2VQM
V46eEcYzP88NInI1JiKJdn2f7/Ko+j2CJNVk5Eeuicm/FndQQlN3l7nzPll/B3+eyDrPRe/shQGu
e5iBHry1xP3nBVZY7o//L7XCDT3JkmaVpgh1GBMGMK+UqibHvfBXDRTbL99tkDdnmHG2z3//TlVc
bnmaPCiT6JTLlE1sk9xaoexM4/hPNk3oUgS2s5xcmQTvjEXnbwMX3/S/uOIVi9mhgBVChj46xHxa
Mxk61g9+SQSO2L0DAjlGB14yVaQO0U1wUiGQm9c++afLt8zuVco8wzZkIzOherypQSsEHWu+9iSz
VKqVE0mULF7yznn3pZ4qe3NlHtEFuACM9uH6jv7sSozy1ZL9hWFP5X/g55uZAnwMRWKto5OXYB0r
b2FQD+zqx3mMDw8U17vjrV8yPij/n1LhTXwDxQojCjVthm6X+l4RQrJbpzTT8GzZeVNbrJ1dNxq2
6/NuddAyMZPVq3kFNaPMArqY5VahK7bGDM1GOZt6Dbm85mPV98Z+LOatMLeVXv5LY+5iHFEhjD22
+6uCLj2WfvgMh52Dh15IeU0fr4f9paNg3f0Cuj47ORGaXBrvsjHM2FGQUDGhcWseWaNTAdYNEHyp
Uv+5oz1C+U5kx6YIALMuqgodnBl+geI+GU5i3mngfvgGPmmYQSynQ4zUV+gpPnfSnAACUhhquwh3
PbpmwXvdFB/5kUwvDUoUjvWqJ1ZigtyWlXhkr+R99y9glkyfpsCZVlADdrL7B91p0K6vAorjTdxa
Hf3j66uIeFjqutV3tIDF74kZxTAfwmo1qJYbVVIR1mCulBUY45aCv/58zSgMzMvqAfF3XlvGWT9S
ebvPWxIzHaW8u/I0fDD5h14BFylFS5wzKHy7Z5Z4V2BfrWngP28ME31a8/nY8EJ1oLgxi/WYP+Y5
9K9ulRIuMk6vi2BChy0UDAjv5W5twYgzKZo+MHz3kd6b65jBDIUDpjijkQ5QoCGDs3Hfg4HWLU6s
+AhpH8WMOW9ar4gkxvCv9Kb8tnu1O6epTVYqXYYDOWEJcLFvfdiZMyUmfgGcqHY6uRVskXhyoZ60
2JWKc0JI4jvsNUNPnOgwKV+EApEWPTuJTzjw5wtHpD90qFMRvkzdqcJ3WaAjZ6kO+2L4PcBIkzhs
S0o4IrOG7j4lvqWShprigbUNPoLighp8JZwzMcfw4ICbdqKmDrG0PMNOFqW5Vr/7X9m1HFoTqpnI
uV0c7xYt3kKesMMHUQsajGCCrtDqvKyky8+0KOG+Uc36TcWqEdM52pRQ7NeaehBcjXcPWgpto3tH
H+SMwiUI5zaX4ZtHGByDImk8Xvc/ri7SbfB+qjqN17+MVCyQR6DmSJI3KHLIctGznIGwRSOGSNwk
xA9+1rtSB8px8+Hhz6OPkBewb8MQrRlO5NjXyPfup2qM/oJO22gLE4EjRQcZ+TekMNYD0GLWBsgH
X6BQnhZy6Q2M5e8v4GfRSgSq5bruK+rWe8BIUa4SZuQtsIxj1wRUAHLTeKOUA9mHqLfC3cA8MbDB
wPNQFVo4k/jRuv+MAWU3pDyy084lpkF0KJRmtlP6Jod8otE9fmIw+eQsrEbyD1j68UQxRLKfWSkP
jb/Y1y9L2PdzKFT7NZ/92qxnJ8M+zqo6iEglAITlhKYXWjTlb4dGMQUsvGaotm0UEzWrY2CbnbKB
NKMXY7zx3jWyy8OHnjY+7FV++m8jXc0aR4hvO2HvX9UPA8w52tMqkkfnlOCeOO3qVTGU5c0j2nYt
tbgvz8w6P+HHNzkIYjiDigbwgFYqXHo9XmOK6n1RKDf0Lw6jRXmeY0jxldNfLH8NBb0wMJftFguX
jGsUkiz0HIkZk057eCZJycuYc5RAFC1Hx87SrwSJ9KMaHbrJ26I56Ndo0IzYTkSy4IuRa8gsPeFd
/Du9w3qGdyj2OiPliVI5Zn6xR9s37rqSOR7xHrqJ9QjCW2EVm5EM4B6NPqcFqfFSJd5ecwwtgBts
e9oJiT387vdRE1sh9AIgYne/lbOrvxC/SfjY7F1JUvtsJZrjmUcgpBVWjER43LVyrABLNLpAUaaa
NqTV63G3iDNvjCBz+DzZjpfEW1A22ris3nZ/ODBGI8XpWc4q/0bANyg6NwUhz+ioJ8jQ3MzB4u2u
QBzWpvvAr4wdHSUC/fmFxjcqIxEZHDBHPFfH7fuMZ2CPhK+l/JsE1wOBxC5sDwrSwqKf7nDvzFC7
MMP/IGUoeP4wjq1g/mXqY0OrmOvB1SxCdx9VHwylmSJA+69cmb5PeRe7vCWoBHRITzYGAn66rW0o
0RcZiy5KOXJnm1vUWlMEYk7HvYR79HI2MHatOiuBXD8dn3dyyGokBUrD/pLZqKNuKXUaGDWurilA
6YmXpEQ91AWYm2fw2Nu0YlzyloHQtbO25F0nwSK9SCXLFvz3eOcoz3PQINzWx/LHp3oRBmtgh+ou
qcU7FFrMb357jY9vYL37hYiZxletCkT27fZsIe3ljwBOKGDkP5+TOXNB+HAUzntQE8hU3dwdGJl/
Z82ZrGbVCsXxtC6oA3hmLEGzOZTDkAd28kaATpMpjPQM/dgY7cU9iXGQ2ogTpuG1EEYul2AmmBGg
ZJ+YT3Tg2RW1aJDQbSrhpMbCP4TdrY7hNNk/wYPzIUoK3E5M/amvxKl57Z21mmBNDyTIG0Jhy7xp
hYV+NQol+Lbts8UOeyoBdn8a7LaD6LfV5jx0QZt64EbhdWbFqwy4ToATCwECJpOQ2GFfnFQOSY7C
PDFuhgNzziDy1rpEJFWunyRNeONTkoLwod5wCmTCEFxBa/bU/I1Hhn9dbfmlO8GqJ6ak178xOB2C
Gn6LqwHd+IWkH+dFTusM3A1mepU1NPb4Na43Xl+snuYztEhNU70Z+22Qh6gqpmx9nimiQN5jeYBV
bfPHaRmlAejOkNzokHfRhGYBe7DSlTNcisFxXlsDiBGqdNdxQCgXBX+K+/TEYhZUnmkqSJ+Cw0sT
lMVK8XjLWl3JQT6daOjpUkkkyZ/LBOp+RDmKcdG7g4//ejFKkdbfhBj8WTHgaFpYpzzKr7QF6XTM
GsolIRRRX+8GTYtH/95DBS4NWLUHUXW4+TG17TcLEXzRq8ghdGPHhJfOl9HFPtFpofzS8qso2Rx4
amL/jO2oJ+foR8Bdx7khciv3+bpRKoQb8KPKx8JCIcx5FdvPDRWzGVWVwDEH1p0d1ilY4FjXndHk
ppojHFNbyNk1Gq1o4X205GOU+3Nj65LrHVpVY1k7NYfJCCC0XxKW2P0ae6aRPH8QzCLBvh3+imuS
sNbpmg+RJiydqW5mUZZObZTO5suyyw5Fln4QTHB9yBnKfmdHiwqdLsiFaHL87NtvtHutKZUIAaF3
84tw0WJZ1+dKoLafgtzzmcuzSoCdzhgdkYbCVvaDqsDFi60YIT/wxpXdWTYl+UlucwKiEIfzQxeN
tdEd/iYAmwxHxbk3exyKybSrZkvhRqahvRS9TyCxkCfIhl8rR/ouNZ87+TLquKMjVqNPQC9c24D/
wrU1AFk6FkQ4sdbkuhtg4V6fkWUTxbUKk6MVRCYEQafkduELjLMBbqAm1kMVlIuwDoOMlXyHvb1u
C4jVyeib6p1astvDaaW3oQqpYft+htfTyOLEUwAHGER8miIxCn8AJp9FgAaHnrk+1orRVKwZXesS
jCmT9lToPhn7WlmYD4Gq23IxurRyTFI4Cwf9jrKhD7o9HhPhJsBCBThHOqdhFwUGDldkmlHZxQXZ
+FmIUnz3EP+QJbcB9r5op1IltrADguFMA3UyIcYcafGKeEFACQDskb12P13GBKOPo6iIa3rWylaD
wXbPlAb0rXYAh9+jSvpvdnBl1Wi7msLQTQKdGaVnc4BOzu/AXqWH0bBtL7xmk2/e8abrx9lJ3xtU
B8UwfIa6eLwTjQA7eHHuZjv02dFQwr73ZYtzhN6QxTCKyU5W/w9IUQMj36xRFG+FcyRWKDW5FWH/
Kh7M2PSTgny54HIBcx3HZBwRfNUsIAav3tvHVW4CmxeA1fKVIQL6OfjiakrDo1mR4iJ+7BLsVsUN
Ze2KUvW819GeFLds5oR6w/MGW5ILnUaTRfsRSss3xY7752fOZ1OsP9CzKYNomY6uvT1doSjjd09Y
l8FPeuNHE8VTreip127LpTFi8iLl8QSISbZB8WKvm98clFo1MNec4lhViQMy8CcCBs2PWih1MinK
d6wKX6lDBzftjIGlK+yHyxM5buuUg/uXZVtL/GyP7eTnmKqxLXPc0mDMxPA4Eaq7O9dc2M3Z6NHx
MNCDBsGdShB5W53ZHICxR3rvM89KrBPlCY2QiBe6Di1ErWvoWyaMYzDTC1F90x5zXymq+9EyKCyU
wEYejvoJbZCRMh6RBXrmG74ukD7640lvoaLMqOoYVXG4VYDa+94XllOTDlqmJePKuhGTNwfLa8Ug
rRBcxj3ePITWCYB1NrhoZ9VVXpyTFt4YcU6ep/FFh7Eh5tEJTU2xxkVJHnxUnJgtPjAFn3JNLbMH
wUZkWr2tjzKkDcG4K9LiWKE8/qVnBY7si44SEkh1LJWfNptNCAenFwft5jG39RNMbOC02b6Xm/Jy
Kb96TkR+sWOPiaDuI4XTtfcNj5LVtbhIWxUHakm3t3OwUqelVA1G0UB03/H6AYEzrzoFGE5u/Fe5
JDiM8Lm+yQRqknou1jTkVUIcOCc0SPdD6BIw3r4368Gq7u2CT413DNRWe53kr2DlCvts9220Ey6X
C2B7gTvK1Vdip55AK+XDWUEPA4E2Jy1V7n6frZFcC8C37eAz9RWOQLjYSYdWYhNQ/c6XOvmtRg1I
QQ8nzg0O/sGiVMjZ+H5tXDp5YPIK2a7MThZyb/c22BO3z9mQ8yXTdNsdElI9PAKQrGobjUXakI2t
J9hHytRI23no7PMm+j153REc7jp2CdMO31ytLkDk/ZCdrzWiziHCNjr8v7dpE6X3Vd8WbKv4eyFi
Fk5qmqVtXzRkGrP7dDfnXgcuEoepcgrVSk3UfGx+hi+IW8KR3hEBxffPGX/JntwzLyRpGeCaGteL
Qgdrashn6jvN0U/iLEoPhI2CH0KjXD1nXr+KN7WpaOI/gkIMCfp4mOR2isTVr2LZYyHSY6xE4POW
+MTJcWFII9PhCbtRE38PtaX+VCSgCKcqkP0ItyYya7xf7pnTr0lzWfaMvBhEe9zp7af6xrrdbI62
W9ormiy5A793wpA/K1T7ZCFREobd0VJJdseEeoZg67ku3gAJETOqc53eiD7BaFmlVdN6tGqOLFf1
xCMTpWmooBseqxEds+OqkoCytWwWI8jjPDJSG6XvMTCBwWPoTYyn5JzxPRpcrgWLwRDL83j5ueym
qgqYCEc+IYIwaae/rOffSTltzT3WQKba1n7aSOVG8UVenM7ILQkTzvbnFSm/XC79+6ryFqijslHy
ifD9Ug73zqgnqIOhWnuQ2jX9udBFNpg22nxLUaTlsiRWzPVdNs5LRBW5TCKork1rMcqOGfWnv7Yx
mMtgIGHClb3odpUXzPN64awdO2ItzO5yHtID2whwXr0+8UClo6lsKaB76CIDxBzOVTjO/9eby/Sn
8L3QM8VtC4d9D73avA2JKpBkTyKGElmVnDxBRZIVWQky1ffJ3MS1D3gGIIZ+4nzp9x/XScaEyxPn
AUUlktgAoKO/E8Q9fyCs6Mk8AgVM66EO2iep8vTGLxqLQlvILsA+0MJTCc3yB2fr5lLarzqa1wx9
gSELVh34Z0AisCIwjzQ/NFrNJMarWL2bdCNSqPG1lZIAdLS+iLUYWwGKwBUszYhlSh++jw+gtRmG
RltB0dvC69IwS0IWAoFsk4EnpXdkcYNy1hz5unvKPuDLrS1sYbDPxLWT0aeIiANjT9etpdJtejzS
qH8RgM1pTkuPxK3w/9SO3v3mxcblIRBQTb958lMJ4oAWtB9r7tUevcpmzteFi1pgqs8F9IOMTBgu
aQe2cba4Iyc5j6jX9IHg5cotYZFA1ZFvndVrV2XDYQzTEdb9njoCp5zQsl3iC44NFHVME8vGdTAh
G43+uegG8By+ERkuJx6OA9QrjrWssrjVYoQmmugwHl9zLGA1NnUf/iyotbaX07ySgRuO0ExUfAGB
qfwSpPGnAQ6p0HA74tqHXkROyyv2ZCuguwZATIOZxIaodtIW9AVyUc6KR0Xg4GBYrR7WH8hhbCHB
8gvwca/3T8BtzIl79cBxPq4KZbZ4oRmC/If9/wLLD03n1TapPHDZ5g/caXC2zP0HyN4zg+Z0knri
Ht+L6ZZlsTjjNbIeabj9mCHbFR3ujp18EBLgSfwAVruybxSddJ89ETx4SIdkLElFvOlbtYb7IRZT
Ulfut2ZLmyNsaxvcHKFfOcMdbA7HqMQUfEdwLix950RBmOyBIrbo7nbW11SH0ptidHh4y14O0eT5
C1pIKoQlfC5bHuViMwnwgRK1Nc11X678eQsKf6JQSCk5sOXl0kzB3974ZidjI9QKgeVi88pHWI2R
Njz1CmjYBqartjpfTRgChwP+/rT7mXNgQMfrX30p4/8PbirN11Lq8BpxoeCgcl5yZ3RgyVAc2nzR
GEpS9Woe6mohhfP3hGGIW1yiBQMMTPVHhdtCLWl6kEOUB42nOP6oawvegp7uwKL34Yhs2C2FY1KI
iB3tOO3v0HcB2TQ9+cLiG10ik/c0Dywx184DFXQUlIk3Ra4mCyihtkBZnho0BNHhUN7LeQNLT87I
8pdLPFDaoGYJ2L3M27/RAPxi5VTxcJeYC9zTx4Ine4UL8lIN7nhXmBM+lNpQqF2NQOAt80WEx7zz
k0gue+2e1qnzpmC/jVmrftATrf/g46badoFmd0A5sJzTNAIG5/BS5kmU+IQO595GZvmJCmtI12BT
UfP3ubuhjW1tQ5FY18lVurMd0rRijCwcl5tT6Kl/uzwLkzahT633mdf442q9FPIJFw14mxUVEI+t
i4zZtjKnduMR8d5Hib9Y6FrIlMK6u9/l1fniX8BSeXEmDvr84FP7rP/pHyqbxpJDitEzVMZugMVF
JRaNXwbyUewrKpOe06w1JYKkjuhPc5GrhFOpIquMN40XjwsTmT1QI3Co4IpISv/3GxWr+tG8f0uw
6ugbEWgQGxSUktymb4JU+V++BdCPW3U21aMxUrKuI1HxuTyJr7hFaGRUdlilsQMn0u2XekQmBMt8
B6J2LXpMlUMRyc8pv/PcX/gf+EuVz2sEBUl4/Dlh8DWCC4q/2+bAdzmVzwu2BhDq3U+StdvMT6y8
KnQDbicRtVH641fC/68h52XDYYkRL2l9fCDGB42b7tadlLEcQYLaNPqlzv+SparQlVgEDM037A35
jOxDNrzKDQ5VmUkxqqwcohWz0KMDi81lBBUX977uweeKDF/fGJgBr1rlRXqUH73VimAgN/aMxnSv
TmZmnS+kxoqVAGW1s8aGtGxHX+sxKkljZJbTfSvAHles3mLlOX3Ah/xux25YwCw2s+ShwEapmBrf
yA2QRyiB8gSItmHPlmApIypriSq5khIsgaxwwvijPM7ZPzCzK5rWMSx15EzpPW8zSJwW30NvEcTv
dPNtyUT/bvpVa23LEw+CbGq2OQXcARfxFIm2ppA4CWjJr43lq3AHr6PI7u1j/JRs/LkjJckO25sG
xxJMI3jSfz7wFb7RqN7zju5nVWu+LDMQAuHw3RybRhQ4oKTtreijsyb53u2msSzegPq67sgTMoBa
kZIHH2jwVp4d5yJntR33434JRoMJSZ29392g/+xu/i2Jm7JVnufeWfJ5RbnahTDEmjaceSPBMvo6
Oa/Ikh2u6JM9RBF30MS7ZIEFBbs5/mKTXFrENliK22+/0RlPtolbmM9kVILzl1Q8sN70sil9ZZxn
7HuHNgIYAb8VozGmKKXS+JpKvul2tJ+QFR3o4ayU0mqllzpC3SKvJ0dLFMZIiyFHrwOvp9XnFO46
p3VYa18FvdXe5JrYgj3Fi0rAUcA6jM2EGlStNLJQS5hnRTiR2Q4IQjMcSlZTssVv4yzXBdms+bq+
hK3HYeE/1fxrjYvohUyomMNzvBFjTqspLrBq5XSObVHjeQqmEbEuDPRndI9qT0jmwjgXPfr/ptAX
Wqf3L5gkpmro5slQy6zt1Y8L+WVGOFXBB73lCILVaRcHWDcxKWYrI2B5Ie13f3+N+hhs42ULeWsb
fOkej6ODSf3MWBfSfv6BiaePIUNlEpn10jjR8AXuReuZ5pDY/eSRfc7Key5LUgGzyDkh7x6lbWLC
Bk1RJPjqEl593Is9U3tXYNX2iQCGepIhxFWLZfnLa0fck0xQ/Eu9UDoFxEtB5GH/ieAGKJ4WddBN
9SgEIEnRyhe6fRcl/9ITfstJO3LFMGhQsskGuR2X2xJebBtWrNrPt/Ux8qwg/IXTg7ii4Yw6z6N1
a0Am09gNuqdnvP4ECsLRoc/pBl7gJBLRPHomsU1QQuXJb7wm9ayKmidWKP4vcqkLYf1h8uAxxIGh
HKOPYs+f3tuh/gkO+swZOfOF6B0OmyRR1pv7WsDDbYAUdpJiwnLM90bm4KKFoTJox8iqH5FF5YIJ
UrIyscsnFpzMzJz7jmBn5bWYz1Fhq4na5sE95/QMrHC5TXvPLlZbsYL/hDy+lchG10WSwypIh2MF
KPUgqqbAoMAg8Z0klZuCSpVGB7QCohx5Z0aikuz7pk9C67pbiz8/RqW0TF36qUFcwPBOrhNsMALx
6EPDDNbltbmvwLRvOJMFwNYZQuHRb5w7PuTvHXRW3M0HyJZNEl1oqofYSjGSAXjED6PQaJkiLvZd
iN1vf/UqI2MR9DOl9GqTQMSZJ1AF1auiZhlfWKk0tVaa4a5jEo2lEKnR8tb8HxRaXa4VodvYpFWv
UyNuCLTJiWmSumAOo4WFsoXtSxPlf1yzxxjYZRHMYbv6573WbVzI+MIem5YOvMkFDcYn0IO1Hs/4
jJgnF/KRh8Ez7c+tM3DANRwC4ogJymJ4ZDrkFpBTQc6spmiguS4RZY/jjXCD81BsxqZuBrx+h5IC
3fLNNa1R1FZKKGfvghn4re+YALz3XZWbR9kwGJIy5WPthlpIJw60/E68sR6UhsikklSuPBnQGgG5
13/coqGZYAJupsz7l3cuPoEYpL+eBF0JnXoQLLGdU/km1/Vpjx6KdkILhIWxgGw9K8SA1AvvPDXq
8jFnK11WwabzX0Ek9tDlGwdb2oN8dsA7Ad+OpKT7ipOKHbNWxoE3eZgQKYnRV2MBVR+5R2x39vQ9
SedoggJ9LeU/zc2wg/rw4tii/wkd5invXD+jTH3UWDDYSjOnBg76pWdsZMeCeEeyqxiIys6tGwmX
IdtBYiaC9hj2IEu0HZy0DF0JealTMU0nepNgVq+McdCBU/scNPEnCoXpaF+sAN/jxfXKi5e3nQ8g
d7rtYYdWGwzchbgUqeBW4xbr/XNhK0TlYwE41vMiwnO9gUF2ZewojbMmOaHF9bQhi6kFh8qK02bq
7iVp+t9AwZmnFvrA7upx4vaOPPecJf/sra2ZpwXhUUNlRpx3Sg4hjCjbTABYj2k+R9CI+3XO6CHi
kqqEXKt8zTN+FlB/yu8+ovrNT7xVnO9MuA5B8uWZlbR7Foh/wC8My4yv9lQtCjIyJY/7EOJhSAQK
Y/LosGlC9Xujx1sJmVId0t2jI7iTTckPPGAKejdudgoQR6I/6+7oMEBjUWA9QqXSij07JqP7ICty
XyIo0uiSLk/IVZfAniULX4PhvlYC9izBoy5eziXFqS/kNqKZrt57EJmWaE48RSGT88xgYbqbvNfH
pKci54Z+KkmDUDmPndaZzquoPaX5k04Bp1+ULl6omShGaCDNGcWFFexDmE8UAEb0mSLHYhO12ckG
+LKyPYj+fTMJD2bUfA6N8N1R0m2Av5Y6uqrpSkMUTxquoRSZkoUnSHSTpSJUeHZ1l91F1hKNbBll
uO/cyP5OKDnHCX9RZx/A19dz1ZoeqwhJWITqZiQKur57Jpq6ahjgFEFTUja/0M0/Nq2tQHO9t2wz
Nj0IkFVqHMeVlR12uREL76MwBUw4clCazJGWDQjLk7UBKA09SNX90O6uGdCRU+0TGxFNcRHrgoIu
hoWJkX3gZyCBschyy5B2Bf7D4D4HipxRNn1xj168MtvKM3RfiMgNFrAgnuBGjGpiwyhQtOyOZVlN
JMWgiOFP5LQ5IUb/X9mjlwgIEsbS1uKGp4CFqCiam1DVVjWszAuj2jyMH7B0g+8YxO7BEjnw41Oc
183lisqN7NhR20+1GJz0T8AksylB3oNfAJ6VTTrGDc7fqveISJXdgO+OvJUmbHuxtJrq4wd/9uXr
OgJMNyNI1pv1qbN7PXZHZ0SlRaLUsj3c6uZD1qM0RjG4st2kda0cDPL+6ct3osMhYpfyfDr/ZgO5
tA2pD3TFF24PxpMr2ETvdpPx69soRrvPEyHSJRlaRvFRUe9fMlbS/1bKRtUaWV5UT5C67GiJoDPg
9HMFC6o06rQLsPr8v/qMDHHg6RT8/xIWAejZr0gEq2FwkKqzm3/MrQj0q9krcb5wIo+b9VC8+p7q
daYt7v1OFNCzIsdS7JUezo/UuLUHNnGEVLs4QGKjybc0iN/1FC2S2npO90cbDoAYsj89VS0b8WbB
h6vRgKSPgbOQc04hZiHBLriRn5w0lyISYxJ1vJwEF5qm0l3IkpF5CkEcAfU0ffq2y6SZOI/ZYx5e
fwNeI/rXNJxa2lzk8yv70ydzkJwtl84SL5pe2xrja3dKQRki49/Vex/tz6W1EdDw1BMqZ5da8WQR
jFb1oInIbQUudS0W+iFWY3uOlKk2u/pTPDqvv+3FwRm9DBc63sxWvQvPcldUn+/OmNWPnk4A1oqj
Sqj/L27z3pwXydzUB3G6M91aBLEBfrmBuMNZoJ8841Hzzf4h37y3mpMGYhMXqvBe7Zv8pEW3E7WX
v/inEJmehmSAl4kewGkP7qXoA281NOScgzrsEwfpiWy9G7jZoF/p09GFEQkd9e4t6w3aGKrsZjnj
7Tt0YgFMziNL3YYdK+dmv4aKSoBwSOA4QngYRX9yMORfVCzdAdsH/qVWfArUXWbLTOGYdJq80qBZ
0yEqHT1HhqCnD76/8ww8sMziOSr2zDxfcYGc8EwnrGL20BbGHKiLEReKIN6OqeBD1LoAGBm22Flt
FTv0iCH0mgvLtFvDHZUTRCCuNUI9AYpUIus1RNLZKCyU1FLEHJkdVXQC5+D2XSOww2D2a1Q873Vt
yt/kK9NWcjbRX8m5PsmV9c/qZW6TcWUgRHYLqiJdVAUVxmNze/Ln7/xZrNEw8RMxVPDDaP5Fh8EQ
7LOaP3XVhy9clGsjKzjNiEU3w82ndrAfx8oJHHGGRX/eZfqAdW52SfoyzzN6J1jF21VT1VNDID+V
C2FzsILHmgmP1Rvm5meki+pApYtgyCLqmsR+OxN/blm7JJjuIvKvQRBcOjRkcZt6hwLXszH7+2sc
a+nycl8phpDLo3kN+hykXAgZVpIVWh7okrrrxRxoONzIR/IFaSQFq2KQv4vwUJdCc+W8VN77PJld
ceSmxtOOhQ98pVyurIdl2bN7sp/189WbQlFgto/UkqZr2h1lulCXD8HhdT9bNLvnb4X9dPdD8ZMR
FKuMQJIAaMP6ADIOUjWYJXpqleVfFEPrBZvYPqLS2xhEx0iEyftTRl7hIDkv4bMNK1Q7az5Ad8G1
wpZLm6cyB7VybPGx5eF+5jTUqk+ywDntEHNwcrEwmwSodX+vBbwIkI32LFn1pCAGSuh7FdJpL9b/
m3/8p1Vyt9wXvyA6WYKfd8auGA3znToq1ee1fMTMUzJ7XOw3GEKcEKclJZZG30d/UoZvDPakENeq
N2nfFKdceOHUxkWQJZ7lxqn+tYiqTyPOC4Yl7VJMc83A3EDHF4MaogmED7SVDHkEQa3sIY5EI1ig
OxoCs1D7CWfnzXEdJQle7dhaK5wXqX39SSTYG5dyJByeRwSQ6Tc76BXKLZgtE07ieCC+IpHzu52u
z5u3A86LTJQYBOy99Gnnnv/vCzWG0JlSf1h8n5kC9qWdEKfYscYQQCBYWn1fGXHEwGs7mjLML8qJ
2YxkqvBhi8jiFVsLK9CUSfoesBUkKjka0IECFa7wsTeT9IHzDYqe5Jujwz3Agqf4QfdUzQ5ZIq7f
tYM2Rzp6zH9oFZnFylpQgGwIrYQO0oLLiU905328o4ZxC238lgv8/YoT7K7Q0jheRf+3LMdebnk1
DQFlDTQvdpz3mPSk24hVQgPGeVKPa17o15Ju4JD2CnTOoHUu5Bd+HliZSwRsEjvUYUsrMWxfkYDN
FuERQ0DHbx7LoDi8ERFm5jtK+eWNyb7IXBQjYWyVh3pysMZoh2L0tl1SmcfD2h0PoeFsgv6dIwgM
2fh8EKT2xo9BH6epXaEXrrxg3skht6Y15OwMq0bds6w54goegpqOI34X8KehPMuJmFl0vq2pDaDv
tbfPup/cG3VvN4vuebGsUN3ENsNw3IUv+b8pQlIqA12GyUZAhGc/nYakKxfcravpFuGD6fSDqRld
3fYrFGNn0Q09JboFDkzDOker7mURidKTjw2M4XQE2vSiu5isw/b0ZN3C+vD2ICcB6/DpSrxGIPbN
R0mnBWU11xOM+GGD+sbl1Z7zFbvWOKFEycDgQhSvTDlRJWRKffCgSj5CZrnglkcetzebv/u6sSQY
YTJH2ucKRfXvydW2zmJrG3A+GoTlDrlbMLuhPnUdN7SWtrhyjGG51DR2qDAgJxUODBV8gZDO58zo
0uSJTkUwBqnE5lfCV1a5ey2MRg6Nb0IttoSOiOoJG7MLZMzjhJ4y5lgToypLKM7g9To9n9ilGl3W
le3eGHumOWzQS75egJeCTYdzOApchwD9p1jr24DLKS6tx+visDr/k/or/wLgnonDSQM5+LV23x3k
UZFlonh8KJ1E7AUdNVXp6MBAWjXWLVKQmNirD9WkLYKkc81Zwzf/8RcKE+XaQRmve6LC0kFJFeQi
CzpDZT/APqv0ddqsb2wmIF/DO2FE/8H+RtmARuzZD5UO4bPWHLO/gHlljfZ+oBmDBwE+Oal2Quag
ejdUgFlJ1Q5LDMXp38Rlvhj/CGFBzPii4N7bMnxfCi8oyu1mpXpttaIAvFXPN6jVY60e1c6+ZjYU
Kvrv2qKE4f5iVMnJ9fGL5ASCPROpGN31QJ+RRId8SrMoqbPmpBstAbuCZ+wWuiAU6nxxvm1bpLNr
KyDp2n6CzA6J+ABVwm+6dePiKAm90qzbmtyx4fjhzb40OVrOIFxPgjSz5LweSQunKxJoeq2FhEk3
a8VNtz+aAt+qFdrHnHiK8i5P5pfDx7DDcdvJF6aUjbfvcn7sLNG+Dnknssl7Yo89XpcVRz0F4XsY
9nTDJFPzT1wouPR9bdgTsxPdsje8yWwLucDMOwIu+Y4VMPmDXUg4ASt1Tmie/prTXTGqQifywUTR
0rslhX6s7dq4cQDrhmIxSfi/RGicAKO1jZdlnZaAqrk+qBYwu5yqaPAzwa56rcPlSt53QZjgWiDZ
AO/8VZztR3zj2CGuy33YSRqb4r72KXQXNS6w0ZTR14WP0eKJ+O+0L2PLHPUPDXqUn/B+hqQDDt3F
9CMXCH/onfZG/KGAaVe0yT2d2YSCQa5eAQioRblOlAKSJFTY+v2R/DtgcstGp9Sf6fFPpTZY5BeV
jkzp2JCzQXVrDk2nLirU1+PUqB62LsRrJaFMH28MqJF201i3truCxTIYQ5d+wURCLiOIRN/yAJ1W
pLRcAaNu5EXd4MtwIhjvZzv3TCx1Qngqo4DRH3pZz10pEOy+X96y6v3oNgI7x1pN0T0sENObRlMi
XuoTKQbmkYWDzXwKomXwhjHTOJx8Zz52y3KQ1TY1e6Ov6GNMSFG5TGf3MSK4KOZKWxYWgTwuAECl
AQpIujTczcfK8DJEFEIxXaO7ygPm6QhPiMt7/xy5NCEm2qzKYDh6K1HVfGfphqHQkk0umXZZE76H
B5dJDbWjCiM1HU/Q280ZqI6IcoCVqoc0jx/6QG1aE9JVvW0q41+sXBTxzOn/IsUQHFgMPC7Jo6SV
ssuuwW+PEv6boL0GoCFWc66jZ/O48VJrgZTG9Mjm9i6jug5jYe6TygAQNlcX0bDMbAfNwOD0MBm5
W4KWybIxIm+l6gMkrrniAC7G9GBB8RUjxgxY/UXhZOI3sD7HTz3FR75OHfx/4Xpd0XrsibcPpnbb
WU7dXdQ6ex1uCTEaiLpmaCrycgsQRsEEQNJlH4ISV0BmhifgGcZzKNTpe45APLzJ/tsWYvznyB45
jjF/6JA+njzcWvYx54tKXLFIrojgYs6rY7yPVADDNr2NEHLQa6UBRDbfxJwKl5pTs1Cdn9J5CL/0
JrJCGOgRSYLFm11psqd52bcT6ZLVAI1qwFaQJ0diEFULBcRSGe5W+Z0ouINT/ZggeKNR31vmqFyG
jc8rWj1vnl8SqxqXvY5M4GBYU9/Jjzp3oEiPb7h8TnGlVbKJ7ssW8PPhggzbKiR0XFJG0YqEsph9
PURWZoFFhTRJrPQhbJBLuahiqXMU9ZTwzCfqyqTHVnWkxlH+KSOS/m0jJeXBzZn3QnE0nrRyju1v
LZ2Kiwl3Of/tfssKdER28RybnCfckHyMBe2inRht4PQ8bOL1vjAGcZYTHjoqRS0bUVh0jhTzu1hZ
X9XVeU25hfC80jW76MrlnkK24XBURITTxAP0lKJVzj71MoA7tg4akhJ+Wb+C6BUqLV91Z/nmEE+c
KIFoFza/5TTTACithBPfjJLtlZxjmYZFf+CyRW2rHJgBXwfR8AujmRzo5NlbrWgS+BoO4EKupsgq
c92fblTa5wtJ8uaeLfP9s7r8Kf2YizXa+OeHZ9xqct/3E7/blEVyGUujJIbxjmGxkHXWUyrAwEzW
5gb6jEbjbmqOtjOL74sTNQAxj+NPkaTCRtXEb9DACFfOMjqu1hlCUt35InWoXqozAU1luneNqjLB
J9vPF2dX0GEl5yCb9v0BE4ZdmTHQF0XtCCxLUhNLv/6/TPM6kZqOjbaxOSmrUuzxUgyrpNCkv3ng
2Dz39uu2YgZEUxu3vsNzzzGVDNHOKv48kBVSpsvRJ53lQ0cPkEF97BEM03lekLTQQyPfcS1J+SwS
BOvB/+SSgzKbGCYa7PNZ3nEjVmtGBYwXCIUQWTMvPDFVta/hzAceKR3o7UfVX78UglRtbFpSATDS
LUdg2c5rkW+zp1jjqYfcK2jqLzDKARUlki46Pi8o470lznCYmYexHPEomSDCFLNz5l+NvlF2Va7e
A6qC38HWOfOnz3tdR++hHbHLYIvr9OB5M5lOsXHq0S/DLH8otmKrPDmLk7C56ZU38vtTmEiWkv0S
BMvKuyytUDPyVpnK/jqFRo/JVmTStJUfZOWG2m/2wzsYyDNzbRiBvOJd2vQHUCarvD/JVf2dhvET
JEBWE1Ou9zHRuKa9UvIfSTuiyZ+WMTlzmv2Pb7WQ4RX175nBFVYLRJj08iIPKrdfAF/PPgWzCpW7
xTkPEJKsa9EbuMKIAMjkJp1OR8lNnA+CQT9JvoV7ShGap6bIJ1D0dYGE2ZBiy3o5vT8hShijUtMj
U6xX+vLyA8ewY71rHC2RCnKIL7bgJv77xUp9eNzWs45Lgk6NUQRwiB5StkNFcWtNgoPSVShvuunn
0jLUYlkcUVVW7I+bbwgerWxyt+U54i1UPD1prvXP3gS0mFvnzFT+2utwVWvx+EDA2m6zIbrzzPDt
a1vX5ms/VBpzfc8+csfE8a1mEu9xdJgjToTRiMYYsCwPQoDSIevJCDje9RvwCEFAAWsm0RA0Cstb
ZSME8x4Mc3OuA0vrXNPGdRaE9G50xHAcmeJnb9l6td95ocktcyuRlUJUQCFo28Eqs3ilN0NSxC6G
zTiRbezWFb8YOGU3JAcCwZ1JgiX4oWSgvTBXLPtPNyTjHovwomJAf/dAV6HIgrLbbs0jvZUVtKEI
BFgrqnxwDUwldY6+8Bumf1My8469Bf50Nsu2gPSbCuUQEfgHHGsTkoRXe3H5fE6R5FSz5DJeGt54
yAjdCub7VTjcCSEvCZ/SSkPbjnlxykYjpVdcRtRZuoTsNo2oQ3uw+6S56riHs6NQkT8410uuWHQy
pf4yDPfVjS5exNUZGtYqmB8PnMcW31nGzsw5ICWBOvvuvD3h1kAdzulP0BGL+vXRnn4qS4ejsHT3
YTzByUgwyCyTucPYM4gyCQ5Q8h2tlrRAyLb7Fw5ug+xCQknj+FRHfvUEN7XdYumDlNRgfGUpUnE+
E2FJhhEpZKLNH0ZUf5BVIRrmzGTZIEy23I5dL5AU8GfiHpI6d5KkCMEZgQwEeAE17bdmPsBjUjyZ
JPwXb4/baM9+ezoKw121iLisf+/d0uzGbv2Ay9ha1UdDLkmkMyyBVWjOPo4jz7G11LpGUalyZQad
evZbMjPclg4UiREtywqNkRIdc+QIGdtgA3tuiJWRRHbMbwgLRrH58fL24/av7A7xdJR985ILtKJt
C2RZsd9v8xR9TLqRSKpaHWvq8DqTmuMtePsqyeMHO+2kYaAPxWuJrFdy+eg+vImRx5m+Tpjfk+He
w/UrmcQsCkZVZMZOS3bYQAMf1g426fa8COf8qeFGv8XV04IpeOHjE0AdamupMPeXQa5V8VZ29Vuj
bD5dQUhZ/vGrd4BKnuT56NEW+lPka7nEWE6WmiQ1wFPE1DOolGUecKSzKIDmJPpQuMKR5gdPVul0
M1uYKwP8My2qJtmj/YAuA+M4UsUdlyJQTyOpOwKdTVR389N+nykWzEyTh27jRkywWZ53vx/7AtZa
f/HmmDOAvcKxFLhdYxP8sVte7sMf7cAXfmh37+l35k36U2Hyy5QcIMNLCjXzHg2T3W1lFmkKu13U
6RQG1Ipb/C4xtjSSxyYjoa3l88534wiThltDPpXH4/LquX3nsQJu0Lq1yl/betYrHcH11SiAufX8
UuvMqEmKYytP5Wcr9ELePibN/5IcOj5EzkingAanKE+BfdcH7uikNxSEVLvJjF7jqoq4S1rEHYf4
uP2WokNlUrScUPIvhMDBlWnBKZTXg/lj8NyQmvL+SSKg/HPpmM8tmXXKIkYG75ZbIDqifr0Kn2k4
IuqC9faJ4HAgiaR/QpSJBWj43RucGE1vbOrlOq3CFQy3gugUgIIiQReJ7egx4D4aM4M6U3kdx5dW
RhmdicJl2IHT93Ad7Sb5xseoT1k8zTqiAr05jbLJIdokp4LfpPQKaalfbpkjyiB+M4jwHqHOOOz4
gy6ZCrPcTelXN1xkXBkSyY6Z3vLkR87nh+hVedJh3ZSIesHX46bHLmzw8xigPg4H1WdOlPgP+G7d
5QaIwWGVXGhy5irUZniOrPqaktRFbSjG03KGUjbR90hWvl8ylzqDg7iG5qDpWQX6PmbTynr4AThT
K05XnzItUwUYP3Yj1Z8LIEFIbyb6cOI4ahbRS779wKe9lqUiG4280OXzNM5bbFh9zqLKKBMiuKzc
uYyNrRO/xpGdVuGIrWg4kpJBIaiswKrhgftT9JmJWmT+/6HYVXSdXlh978EE9Yi1XGpjLbmg2OnM
gSZ64gWecmCbQVXvRoWN6Aeoq21QUcjDlg0wKu8YnJ1xxsZ5LwcvZ8usI9/PUg1cHLioFMHpaGiP
jMps7nXsFyNwP04p6rtGsoIa6oJWa30p2MGgPrPqjlNabAbCIrZ2HVok4QrkXnQR/rlSwi414Nsy
5vJ5ffOg7nsAcrZoAU2ZIpxcqARL4tVKmV3Ulu/10KXUFw9OQavg4q7L5qjSAsVwvPCXbFin56jI
Abosz70Cu/h2ueLLkdD23h3cXho0q6rdgBWZZzGrM+q4NH04I/KLoGSN2n+DLSnKLGn4HcQukAiG
jfeJJig2AT8eqoHoDxG4ZBDijJcSM8lZFqGxYJGeymSrjL1r3SgkQ1eEU8+4JtLaGFypsROjWbjF
tA1xq4JrX+OCMxYLnrjyD/ONs3Rm9WdSmeM7cW/ssX+cJUaHJ8JPtJQZiY9Dv4cQSEueN9StFKVg
Vy5lKneh3Y2668Nuhw4ppi9hVSqcHH2N30sPC5tWKa/Bu7xS5gYRhywaVgbVd+4hOs63Xo8vPLlI
2aw4XazRojjGtzMdZqoE9G6KdMzi+YEGgyrIzFGC55T85+ybRBlKKktX5nu+6G4aF3hKb/4iot30
cpMN+/Cvm22ao8gF7CiBcypFAIB0RSFkhhA34YP9c0UapXdOeDfadVjSnEDTQI03aWk8sDQJ518B
Sxa7BR1OSl4bx7D5LdkyyvxW2hgX4DsubElFGdgkVPbag+U7VOaUcgaXctRI2QnI8nrhWFmRUQpQ
FB/gMuNOO1YK/myoS6AOU93/TY7WHS9MnKrhmENbImVP2RfVJqplTWlfDLAB3az5mmzdpYekQ8a8
AjqNmNDM2EYRGCNQIY2Paw/3dYaodtQMgG9pDxMplLTRO4FqGaKSQ8PofGsBAWmJQJwE67AI596N
ynneCttLdT2dbuq7gFfuGUzKNS8mGpUxNdT7Sa0FZns68Nw4V9W1HUysY1FxsQiqvij9qGuIEAhn
RJFkq73GUba5uyaegOXY2hcmWJwrPG8x3f6l57QEU05IbIPerEK+tmzYhAvebA2o0bYVox0zYI5N
2sGNCmXS8A/uCCBoQaXh4dM5B/9ifHoI1u3D+NsVfFjHGcskvwsY4lSCGHAbgda0hJK0CnF0mi2O
UE1L85r49KwtMtp/A/G2V/IH6inwXB8HX7l0fMoIfDLDJh9AWiXNSMGsf3td70czbeTTNNxlem30
PoAby7+7J4q5uJc+mWtxYqJTJKPvmAtj2TsRk1FAns3Zq2qJUPIraOeS8CYgcAIVnpUstUIKQO/i
m6EIjjTWHvkwYMJG0avQYFbo8Ko9QksgY30S9DBtn18hKSkm5/KNrzAJ3HkNqyAxsOvEoyltTwER
gCraxVdNDQGpGg/rIThqXJW7cO8OBkHa2ydx/pc2IxpxnwxuXkppXGpf9y7E8rebOWryEIs/NZ+W
towFHDvqcWbHdx9U8GDfbnfOer1vAfy2eanPDBOF/GuxIqtZoOVgIOOK36lFdsYQJxB0+AxP182E
8tRsKXVXwJnQtlnRRkavKjxCCOIT/WlSx00FT9tizv/WK5mPPensXU3pOlyUazg2gaavFPfI47Er
l+J9sBIziA9MISifeRxdoMCJgfg23/8BhE5Rfx/g9F0W8boLa+a9a8fnzkKNR72xkJZ0YsklQf/W
3T+jrmN4wgRVgAd0L22Fcmjl0BkwVjgo//su4uN4oD/A5J2281+CFd5FNM7fsEh5tJ7bH647nM2F
Y+r0Jnrn0KBR7m7HIfYLW23UOQt8uTqdL3NcIvK9xhCbq3jUvgSPNY0rIK7KuoLuMFAS65zrkBSZ
ZEluy8RspI13pzbMmFLZosWsKusiKB8Omb2rwXAjSNN/1TlB9W4HrlDxNVCBgSM2CTsioGiddtnp
trUqTVXw5KP/I2yb7J7Y4ygWkT5QHxSJKyBgYNZ5AQIsQoq35CWkrXY49TMdxTJ/EREI0VwMyoG6
qmDPKO6/CxI0MMi7dN7dw6tfwlXNWEd4KIjn10QBYlJdCLIVgv52hDWglhKL+lReSs6fSPQ5ds/o
X6zXuIZPB+Mf7t3BK0png5tjDkqc+YkW9L3H6kUWGNdADi8HyYZlCcJq4ymavQ8LfUtaj53cUUW9
0npTOU49wtVqRSZPXTbiTrtqmdEWmllJF/GyP5mFiQHRsI6HHvN/R7ZkEtc+M93dZLO2gsnciCo3
5wdDcWFj1eViciJFw+s4J+bPG4+eZ8pQBGWbELQ/Uyug1KLHBqLYUGy9I34blz35vI0tXFCKs0eW
ypQQ94l1dkaNCxVBLrOZ51aXKYjUd3ME9gNlKQTWH+a/N+l+B+W28xk28AXRb3fuZMDmh77Ftyoi
wfyb1SFm+6fJcjeOwpkdfrYmcyWDo55PWnzL19uerCmvzepGtTB7D98WuenPltWNTS6gFGuo+NKO
3dd4VHPsxnMSOZ1aFAJk4PVJjDku1I9t+6LOUe55McqgMIaUVWqBmQpOkY3avkrkceC4JsGyr8Cp
0MuAIn1+mpUPOK2zjlMJPOFidYLQ/HBIu1TxcUS+o6YsO96ZlLkhVOAd++Va9K4SRUPwqZXr34KH
dIUdqjYLh3zK58MCmlXhuiQy39+TdbiNxmyIqwgiCbfFJiO8/xfGEfmbpkNa2nW9m/6s7Eycc5gM
9OHogZDJNcbzJ/JrjjxWhhc4K3hYs9mfg8HsFS+6jKOM4Qkg6ETpESiGpym0D5itJJFPz0A9VWe2
VAtJYakwi6PqFk+5sSlIXHwFpQKL2Nx2UWnGsLMx2lPJGGRF+Bx3+iayGiYvJyaY6P926RdUTqV5
3S5MGkOm/78TG+8pp0zYN9s3HyfJubrVwTzgW3sLQ6Rg6YeFvF9CejS7gp0FytcPQhBibHPt+AoQ
64jkl8rYRGu3qepQTBld5ywj6I0a5W11rW5NtA1bbyFox3TCOrhKvxgVX0ZS1lAAVVikvyuksSDO
nAuBjYpdVmQM+UmpqhLE9jfgJ9yWNRqHaQRfpyxuOWmUQMd7oAN3/GVQdAPGgTdFGWRN7lQ8z5qP
+xYrWi09ciGeUNeYi+f7gfdIfKHuepRyDifhdL8fwwIxDKYpcqFIzlmspsh/I2h0SQA6xPOpevli
mFhS/8UxjbHm5INQkwzJ0PHbB5GpHFgdLDPmYvvtyWeqkwBzMMMEl9vaaaBFH0DOrlBJ0Qa59GBT
3KvcLWi0CsrVH7gK7y7pc0/IBt6YclBhAavN9MABP/tN/E5Uz8Dc/lV8lhi0G6Tizbont6ChJlLz
iGzXd+MsHwAknJe+DoyTJCo0zS+iUvXrvZVkrRJmPeTuvyqQ5t1DLqedGQ9jyhzWv0pT0eSBmPWq
Lzkv4vdO1ZZcJJoaDN44yIqRIfXoiAGGdl7dCzO9V30QWVbaHRWXcVs32BQJam3qGZbf8m4xwigL
35Jd8GkJmsgVcZgCitWJtvFGhaQiUG4Oby14jzVZitKxupt1Y0LXEptsz4V0DbHnXdaJkiNwloV5
28OUDst7FpCJnp/PwEqtY4//e0hQGwq+6ed77FX1fpIYkOhcovErJKUjGE24tceLSiOtGxQPEvDT
b8A+XA66MVzjtpT090NbO80XZM4tAOUptWEiu1KSraJKpmmMRqGjj+ro7qO4dryxA3rNL4svjO9T
0NbNeTdjKJRxzIrgRQJ0kIW23m973lsig1pKNlWCA6iJ7DmoB5+UgDNWLTB0AczrrAm1uNFCX4+4
sJGN5gcgcx00Me7CRaWI979oc9vHMwT9Vca6GpOl9s5Mne4XgouVSBgTzTItGiwDi5AnHy5XPO7R
sOc/Snd3pf1YEXzFRdYkklrMbiIF3NtqmoivioN+hfsk3ExReIONC/6FJ+hj+k3iAlQ4F0tohNCV
LLnhHYWVOo/lCHnTreW6whIAflfevIao4zdVtNfZHtvvYyNARBIYoPHU8Yb4MGAS7+VulCvxXZB+
mqGk2lPvUi0J3DstoiFbeCYLNthkhnG/wDTIPwCsQuwwnswa1gnPi3PEP19cM49kFVvRNvcW50qp
g3On/6CKRfGmv94b+igldq/Umai1aMXyAlkiI5Cf4APPWmKKXmgNyCQC7RqeP9xSEz6Lxb3iRXlx
TTyr2DxyHwc4TMKYXo/fOJDFob9jdZuplPwsQAp1GgzuJ9XnFv3YdTHIVk+2VmprqobbglySUY0S
vFEykqd4nufs3l69RKmv5MAjq2aNzHsDAggz0hCtnCFvlUw3OhXY9JO5yeedkhkRwI6JOUuTD3/X
1CGQbYAWh1IbquE2XX6F4mXTBBvSuVcqlISCvi5uadAx6maHsqpL/nOoinSFOE5B9qPOvZXa60iO
9X+owLRNG3AB6+4/W2MB4t6x7EzGOYNQ7kNPdaBkLJh8dYSJR6FNH/pqaS7QA7h6LB5rQOqCoF9K
3BYXbEQzNavs5VcaZrUV+zs3iBHrBG4ponNUlFbGFiYxf5JgJU5P+vEqEpCjSSVTUspV3+3EAfLj
wUITSrj93COVZOAC0MELKhewi3mwITKxNddMeXBG3SRTKu+KPvYC7Qn+FJaeMfI4XS1WPKY806ZO
l14Kk23fM30KpK4uzrsw+r55e/nLwuKbED+VY7osO8ERTtc//ksKvnaEHeaPn0tSWXmmNwS6tb3H
GBaq5ASXcaedZBhvClED7ldrlzA2UwJPPBR86dCt9rg8hY8kXYmS9jbhtDw6p0cb0+GrGjrnkBJB
LHSbr0Dg/sfFGm24gSfq5kElJWuGGxqSnIFfUBGhJpnU5QQ1iRggZ1r9xjR3S65NW3S7iF5Ek2ln
mkRD5M1k6Tn8qfJPSgbA5DzTg2fAzxwc11BuQ4GcFpzJaIdJsJOq9SNXAu4wM86F+hLrpGSYvJAT
b3sEFS8/fRTaeHJO+nppKeeAqoPemyNt5nzZ6TCHuzgHLLL4MUz3sPMQBQwpQRnlDOKfwe7x6MTm
JJVmEPH7bzO1bLhzJ8pac3oSfyQA74oKvElra4JWJhhM+TS1cHsV/ttqJ34wl9Z33YO6da46y7te
Q2xFGnl0LXz++/a2eumuot/dTYCmDMD4GHXvLS+84bhq2zM+I4EH+l414BgXymdggrAZpejKvPPz
sF0JC66IZnXnU8ZuiwfWrojaeV1n2uB/rlco5nsONwrYy7iWoYVi0kRg9d/ncq1LpUVPwSeL+t0r
6IJKMi8K8YO3Cs790GcclufAju6fI5e2zEghyR9XY4wGz3WXyz4lt9uGmVAxlHDn/liiUr5lY0+f
J2y8vY8YeDby+gk3O7hGm0f6aOlf91BeQEWxQi/CMp1R8BeVwI3rKvgTjswQLzrbxpFRHB1j9IHj
qbMX2lfXs79nOBnupf5FXurkP/mbpJ5y6zQH8gpfIv6EFZ7Cpm1vVz5svOHJOZXaVM8NyalZEMOb
ZdoIBGVqh8iqORdhj765a316Ftx3MkTHIY3ePndHXnm5KSdVoAjj8fFfQbKqMUtrqAIaU0+LUwyx
c/EdsiH0e7EbwyI2CQ1ezECoZghhIWQMhzJscqj9wEq0q9m+jRayeEjwJEuK+Kpq3O0zqCbKT9Cu
uiQNafTeVgsHiW2cs0epo+TYbKqo6T2khLXYtkF5jUrvNW2jB8GHGsASqPJdYmjLV03L9VP7Lv5c
z2/CpauuyWbG40ard1sRj4pqm7dQ9MSJ/O6IJ4HszvFORFLfgMwgAFxnkoAfBBkr3QnUPMhQxAQS
TIXR18UcTdnioAOh5U7W8hq16wkaJzVQ3hGLgBxqJs13b+nPjG+Lpyg/CydSInmcFwp8KxRPvJ8X
Fq5fvEMTDjf9hfeOXn0Mi1h1YzScuM2hqgT1f2XM2qzXZjTFdKfF3/icDeHulcAByAPHcCCRqfTA
/T5c2k5Gjj7nbcJ4c0tdQM/BwP+etkB319wKhe9kK5x2X4cAwN7JjDamSvfuboUFXS0JiTHV04tq
pMRK16flB5Bx8t0E28WyoLTDx1aHB24ISFVx97y4N9b8NqWiKcNQIW78Q9XOMnult1MTqSCd79NI
+4vXxhWLXGjb7/lniUDa1dnwn4qHJkiVyjTNHl84mB6smEBmpQzcXWmPpExScinLo93qHCOF1bdW
R0s3OFdgZ/1F8LzIvY3f9zbp5jCznliHFjeAgQpkg660cxievzaGww3GTYM4deHWNejY1tqyVHhe
WUXIF9cdE4ctZ1ILC21OXEIPWXf6lK+/TjrP+TCuRKk5D2WVGvt0fVutqag+ODj9oDNe3GlIjUiQ
fdmgOuNvjkZF/WRs92NSDOJBhBL9zP9Ui+9Fb8iR2txO7BdlD8Pp/yn97oWWe/GpeSFhvn+zRAja
lsuAX8FU72O9jzZAM45BdbKz8rlYJMN2oExN/HY4Wg0XqAPFFuhgpiPYyEDl2PhT+mWhgBUaDgrS
9goRjIkERRuYmVrq54XJBJkLwbFeAVABMxP0Fb+wU16AzJHZvdyNNCbCSVJwnzKdNb/OfOYIGqhX
x/tp7FKlo0+NGsSitP2TPyRfo2gJ4yA0aPenhgUbu0YSLiKZws0w299YEP0b7SkIwzYtFR8OefGN
vC/GqvG8kZOd2K4x+VauqojXRdSsflprf7o0jfcNxWpvK7awOHFK4QjPv/MOl7hs/GPawlcjg4uf
JlNlf8MS9wgU35f08RFHC3D6vNqNnc7wXLnJqBC2JmigGmE6JvuYUbqRelf3NVqOd7/VSYawpGFK
j+EA94SpX277TgZCTfWVeYvyYfU0GI9EwAvYMiKF+tnc1raBZ7beum95hEYDAQiqbMvwITgJfM7M
O6HS0JTUNg9Q3uSnEER5Qb2oDKxTh4UZvZ1kHEfFxIlABh8KfUeoxVGV2zSWgKGXHfRTkeNVXWR1
+DDlo7TKbeU3NAxoyuEEGD071SVqVR09JLgrKiNt8pfm1FXf3vkz+gwekDajktjjRKO/jZIl1o5a
5tgNJPq1AxrervDJo09Q1q3nQNSsif+dr6D6sqaKxkHyRdshtPM3fRltm/1+vl8p/5d5k6lTccGz
t5g7zvD2Mw4CCW1SvhJGiUFFGuu472ut62pD40xVKCYcKCm8xHogugiLqJLSLcUtHOb3SioRC9cp
VryvsayHj+fgmITQirb1uOaJLuXW2GFdXTx6BJ8OP0V5EOFmZohuLkut1cqLVSUTWW95qKltb1jP
erES0VKE0ZTnzxig8wXbjmijLoPtLeX0544RLw4O6bvTiWjJFpGZD5IDJwZL2p9t/0HfcgDMA2X+
b413hOHMFaSCdnMiP7aPIjjPHkPSshoXLyEruQKc95BSNUIMkrIX7CFC3bgo1QVsmbuAdOY+KfNa
6e7ihFLlAAl8RNvz7aVGd0Buiv6lavefPJpa8Y7qqw3BNdvllMj7GdxoqrMuQk6zw5eXiZcwidaF
+0aTsdAhn364m5WNj7qPXjne0h1yAqE0OHD/VhmkGjD6PQ6BvRUJ9e8d7uRm4TvOCHD0Mq+jw/lJ
hb+njf9RerWVPwxfhcoHze5WZWP+V4f9PU7ZHicUAgqS6nPphpbqDQlXUAOzc2UgHan5koi8sD5o
2loPXOh9vEnj5UtBvjs6LMDZLmBAQWUs3xFEBiW0wWHfPLX3ZIPinfbgDeLoAMwcVOQUYz4Dvjdu
XGIKhHmhMMNVXjamOJZ1ZgbJkD0HNjjF7fLTqhGU6GSuJwFyU7TiqtkF6+naNU+m2Zq+rGtUK0gu
j4V9ekENw1fA/Y+BRs8ubtq/EzNBHwTRGcGe3LN3X3vgQ6Td4rLam3iGXtK1w1rtuOxpF7HBVrGE
4xvNs07ktDvwHeHeXQCUKQCR290cAoFiIGmf9rTcr34W4LBEp7UUZ23uirlfbGYm7YSlj0BCsHlu
2qTQY7Ne6dEyexWiJQrCDQJVsi5yoXVDyAPC5H0gpes0sSjuNb+yABbRi+BKlmZJtFsUJuFRCJxU
MvRqtBGPWu9d2si2cbIisItjrGSbRWNEyYrxki5O5jVPq2VGVQnoo4KtFd2wxRdO9QyprEVslenN
kfnlZfIv/nrFTEShgcBQ+x6ZiB42w4cZx5RigDFQjglB5P66ugOuAQ8uZyWNxz4zhKjOezcZl6N4
WdM/KuTe2kmsYkOcQ4Ircf6kYT40lv3k+KrFctGxgxc74FovdKCSKQGdcpA9acuO3CrtPFZgy+cA
fWAIIZhp6oAYbTsdzEfe1csYkb8CnsnEmdGDGodk5rU8Ts5SWQ4c5IkESKCQQFcd7+Xt0mqIiI1e
eHIFW8VQBTU+DZ3MDkGhSl2IHHO3MxzaaDlIWty9gbcH00YDE0FxrEpbN/9d3utCAHZQzD1kDVhN
6Xtgyr5yy+gg/mdMlSEZKIhtMJTlVyVx8wzIwVYpeKcn0CxH/tai3A9nCvllxnRjfqTO43qZgvF3
KIw81YrMk8W0bQbNHT3yNJ6tdGXtKqmYa/D3OnuL4T4+204Fqm2qKA5rigPdXDSDFfLqnbHIz1Yx
15hkTHHZ86VDThrwLpWskvbScWwB1ZcCdknfJ1UTz02Guw0r0iXd8ltQAW2TUipKlkjAx7F31MG+
jfN1ZyJtCm1F8P8O1PuTAVob8KbK6duEldX5GFh+9wmWp8NEm0TUln/aEYR7Xtej501AKxVtnwCY
oXodv3RAUtGkxRg/K3a3Q7nSjejwQ6AcwZD3/P7naiw/rLq2uN4IHHyjkV83rpVv0oZuvyPX0mBR
qWh1/O71xDqQuZFa35iWm3FbvhMG7O2X5uwvBhxvZLJn336aj80YA2MDVvV/2L1pWV7X6zh5ep+U
xs0UirVL8PJA88t9++rKNmdu5OjNG0JxxA8k+qRBh/YmE3wi4R+4YkggkO38GHtGrNSu6noXHipS
1YG1KQr9K51ocH5W0ebY9GjK4XRb7DnKaHJ9BPRjrk/Iv7gN5XflLGlFWgY4PG2pAeTF5D1Hjsi3
YGOr/SQYzUdtKbZQ6EIFSwS1ZRGxHuBJKJSmAyujmiiWQy7NcZ+y31ZwfNMhMlSOs7FSabTzCjvn
JLOV968tWyYOU9AWGdP1AHgpSOW86zbQdzqKF2/hr9Al7Siis9cVm9D2reP+UBQEMZdktvkYjhBH
QqGwZoR+/D5bNZoGFZ6Mw0qKMRCOlmw+4dgw8YlrfFb5jDRcwVMFxwhitpnbcjnzcCOKRTN6sznF
h69S9NvWOfAQ+3neYW3OWTNXoFD7RQV/Nn0bVcffKFyWUehM4g+VujyVf8+T35wF/uksEa08Xoja
EuMh9ri5R+0NqaJ2gJIx4YalZst/ad/BFvCFJv2Zp/vGKi3VqwO4qpdqkt5BiGRXvbzBXd8WvpCB
/d9UMVSSzcKp+PKJuxhuSiBHlBA4a8+KPBxcNUxIX8JN/AvsLhFzxmxWkt5XnnDS3k/zE3NMXUY5
g1wx+KXrzMlvz/R24aQ8DVT/aHD0uXWwjM0Jrihu/BCpHEP++IqVKV6BHHnxB6qkgnBMWNyPksJt
3kNOUIvVGLXOuZh2lUOX4tbKyrQfFexWJf3+DAC6mxzYPN16v97qVeEvXiMlCzNk3V+F4QLwnPva
xhoylxLu+2c9JELVdxVylCl+N+VmvhiP58q6IRMRZhGpVsLw1DkUUPwAHT7N0eYKMBJT//1mqQ8R
8Aok1Z5Cz0DVhW7SV1aVZbW2vQAwKzLsPlqUBh7Vz9U+zIkSvD/eR/P0j5JM05wJnOPaAd+vxw3W
0xI/d25WD7vfPZpcBfAk6tACBYwZryxnRc2h0eaSKEHEinKMoPx7OdeGC8rSt+hssxjXlSVh4BV3
RfwK6/QVG7hfEReF6XEioOQBO7ZXNqcvcDa1Ran85pmWrQMkvXdRk1NbJSebxXWNl4ooUULsP+Zj
djg5bDKb2DHUE35g7lkln3Y7igDAeqHWX7eHD9UvETekF4OiKEGs3FIuso5l3gJMfTO4l6aAtvVY
9b5gaC8nG8CTS/twdA+72AVGMMIXQ1KKg7NMYHw6CNSBTDMkdh8yIYbCFQ0B8hPcGywXu+llS2/d
N7wIpPQxbq1V7ULfzq80dRiCtMYUgTCgQNP4odkOnPBiMNJfZgRByw5Hp/Uku7A6Zhed/xytzjC5
R2IuvAACM5ypxdnDkRA+ueHqqygLzteWYxiHXQcQL2NhCEaMBIREN4PzrO3knhS/yEJLXldxquqs
tr/7JW6wQ85KjxwOVe98HgMO+2Aj9gOvBBnETXxLIRAULEnxhQSKqQ9Ja4z6fWvtuJOLUg1JG+8U
6y6ooobatkOaVIW+0Bzgrb05cla9b3OxyHXcfw9HeThW6V/pDgXgKvLp41mOfXDRi7v7VfPy2Lhj
T783xCnv28SJyVRbrKfjEOL1r1M6vh2gDE94IFCVex3hOQjg59K126pCqTVDGV+HcHfHJnHKddAW
SV/ZNYLmEe21hHyQXiiG5KgbfrXhy+vglP2mMDZuQiPJ4sUolkBOSFFOrFRE8r//OoAbb4Y89JBo
Mkq6O6lwNL90mjrphivhmK4hCB64xRxa8K6c6ykywMo4QgGEtcHBnqq8HEI73nVWFjW4RIM9JKPp
FWg4rkgPBiAjH5XawT16DvKAOgMnWm18Nas2MMMmcaEVOtJaoGr8d5VMvDpIRWTC4XtyfsMeMvog
8KR2gY5+7pVdzPXd03oQzU6ylYFD3JOueh8Wlh/H6W+EbtOrh5TQw406ek+fdDy8Zp4mDtcUvWoE
yzbg0NutQth/J/k46OEjANaACwaC4TeXHtPg8rIlRo4D3zgUPLNHGTl63OQ14cfsZDDm7kceRCbK
/C/pnj7ja+WJXmcHrSHAompxHlpQdWsn/esiTeAKLE2vseSTf3zDsnczqe3AOsoVYkD5jIQl5nzH
dSN6QkYjSnx1wHtQJB3pft9WAugA3UCUixbtvV5nyu5dzMCK9l8Ix9+cGkwnH/7wjkyJhpxwPBUF
uQgxFGP6EYunNSUY5C3CmVXhJi2xrEjPNfRD7fM+nBW0P2kUUWjPCBj7Few8QyTzKv/Poyx2xyfa
dRjvu8v4eRsmT2/2zuLk0tUqc/p2b6poHs9RR6bejd0nW1CyRLitbfRpzcfjIfau2tWAMMWKgmEv
aau1bMB/GetyUHYt6xmU/NPhmQwbHVrOqasbqVGYefPujaUUq90lmBy/yrB9yziVFJwCNn2V5dBq
v9xfR5sXvg+Hoe0A5VOh91Itw0srQFX0m3ScrIFHBGOP5QknWeekJac757wbvgskaaCF/J6nfNhc
WU00d3JdILGTV200d4x7sNYzYjYk+zj1Q51mNyR1t5WKzmks6jEJQN3Wd+b4ZlLMdcgNOoNNkIPc
r/Nh5Q7CeuY5vaxyMFMTrqF14bC1vcxyh9z05eO+wNZhMMdayQ3fA8MA0Ch2PPRCyQa4QCJQNHo5
h1gdNyyiCk7ucSSlSCbKNQ+XP0uXHOLyEWB1bHV3TuEXoogsJot6QWfh330ocAXCYSLNwhzBJjqI
Z5Cs/h2aGhXvR4rZGDXcD3u3/6CHNyvQIwx6TwR0TF3rpDuuf12iKO9TqaFPGOg/VX2b3hUN99aX
lxaKyq/GOLRSgHb+SuFOS1HgQ7B3AggJOoxhc5N4QZlX5OVpHQhtBhKBrtS9CIls2KQJANJVjyM6
2jaASSz4/lcZs2XzMMv+87DNM4XJAksUsnmBsLhFfz9jpRJ/iE/Em+vs3QrVMpyQcxWujHsRlRGL
BjfDOel33BuEF4R6G+4mpJahD9GTcmgxTsJ1Yjg/QZMJjEq6Zic1M7tpEJJmZHQeYILJXXZGrxmN
y8StEZ+R7BZ8QhLAwlJ3BWLGhoHqacq6YvNzbPvUSRud65H9tvQJcDKhpdv086Expiea1rxHWwzO
e7qRCL7c28lwlW7n4HzovSBNxrDQRbh2ZLPW0IXctOnBfV+1pS5XpbnHC9bVKtUgRT7j0ABDDcyc
Gvf2h8ainPt4ZHwsQ0hpLBVLKl2dSh11mHOx0zTdA8zcmbICrFJXlVxNIoeiIoqTJoZ/ESYLEp6W
uAFNKQRXwFuM3W7/BYQW9SaxbMzD+bUeg10wruH9KemBew+/vQ62qq6d+Zd+QGi3Rsu2HwaYKAbi
h2ARuKDRfEYVtXQxlTxYdyz4FVx8yGffukmu6N2UsUnvSGI9HvVk9MT32r0e8iYMldQI9ud+YB5I
P9lG/mYLk3Pkl5Bc2kkX1mYml2XWPtKu17Jyk8oRW+oBVhRqF6e7XjV7H3RqgrhbX3uDAPzHO/9p
Dk4xZiR0Ul0ENeicuGAt8jfuPJzm2BiKxwo0DEgrlYNWo4ltsuyh+7F7nCJRRCOI+68/CfJnk6Tm
iP/B6K/408nhp21iFqh1jhG42rydliewmKAFMgcEepDNpv9fFwXK/6iIxE+yPAnkskX+QNbfddbw
SHQLVEtfmnmxBvxUow7w0pRv0MdgkE7GVZOvIVTmv9kHpCu+RkevygQNnKGC2ojvxb2PwZfHlipy
gF+NBQltHHgcDUw7HjJWVunPnARpU7pwvXeEEnfx64jTV+d9cDp9/2arqZ1ngJ7ax2tl/4Kk7t1b
Axj3VaVx0dvPIjnrjqbten/GqFbe0aMBx7uiEHnyUbZYxuGRzaHUPOZZSP7HHDdYkx8m8gPXutL/
qLTIVsmNOu/UxojnBbwNJSzRjUcyZII66oMppia++0UWEaqHOB2j2xmrjS/AeVVLrEbTHSWfs8/x
XcUMqB7TIfROdPZbfOl9shJ2kx8YEHimrZUcJBzzJ5feb7r4wCoViY9NxDiSaJAIGBe4DD+0EFbK
SlDoA3rhYsnG5pSEF8LuZsoY6GyLovn6FiuEEH8ZwjpZHTMgGQ28J31W1xE5jJ4ZbA0W1DLbYqOH
NGqUvpESL7fz8nj0ZfAA+gDk+t7gnKxazKKASyJgwcSgl7vOz74LBKE1jRPhJ0dZxIHoaQ04nvTm
WUpg4xG11wwJkRsN88+4jpgg57lf9CRGpH2kE1olcyxE/hyYwWNhL2EEuMfXtWeBVfgT0mwSPxBd
BFTmBqPQPKUmH22Pgo5Gl4VjILJU9SHmGTwIgemTrnmsXIOLIlSpK+bUxlnmRvZ5UhjgbqZ1Bm67
tYAUho0hzlKmbVQvQmElkL6WfRQcd+kJQ2cNQ+xrkUjwwxEBuzqaZGuaQbh1OmTroWpOTbvuzCac
ZhQQoazJOxA/gGxr0bGaSzB6OLT/qgzHH0Cp+e6tN7r5MyVcjKj7TuTUBJmKAxONm1IXaQ/N2UE2
K7vXB3SP3z+/rnBV4ggblbyrlo3WoapdSzXmRa8m1T1hk2/g7MzrdOHoiX9IojlP54Ejru3sket2
gbqGjdvHhjj7OxF2Mfh/mTYhuMaBPeuhJxcOekWuEIypO28W9yHhSd8qfy7MkcvCeNnLOyx7LnGB
Vvp4r1zxrcjtd/Hj76Xb5dr7koxodoeg5HTmqihHB/QOnEHgs5lNZYTLcHuwNEZG/6ZfIhjJe85e
ox0AXwfFG8Nxvpyzt5FahEj4fIr1LGPOOLlGBg/8LNior2C84yY+yBY27KQUXiVEdD/pXbDOzuHq
xGU1V/t9eXNmXs8xttCWRW2dvPhahjDBCQFl4znuc5AlDHqpg3sLP0pjFntFkvkMpHv8/47+1agx
3pZDhIi+ho4IUegnXIcZH7yBwO4DNRGUpPt7LT+lXx4wfivzjFyjrZVojCPaqXzumQhC/kWC50Lo
/gpCmizIZBWyRO5JwRyY8DtcHKd8Pow6HUhsobcnmWj+z2FbFJnT8PaDZIlgEEENlFsvW9ghsNxA
aWST3GAIcWNOqFAh9z7S5+Llz07aRfsitiDW9ssizknrNl6JiuMHIJbGfUyc1JVU1q6yCZb2VqUQ
K/dDmnBVtKzc9PZJjrYAIQiUgL/azNx1vygahggyn1ZTtLhhUY9MlI8u4Wiuvcua7Sus8fE5p4Et
UBOiXjmQNqkMp+ywOaG+TMqzFIfkXBgJ0KumXWwV/8DELmZaB9U3QCEqoPDBz+XONHZ+2wgyJNxF
Q6j0VSZZHgzasTDLc18SmXAd+L0FIe1HIjI30CUlEMMa+qwQpt1zswI566NS3S8xPDhQEfwf3bIv
aMJnDOFZ9jitSrXM+YKbSPSKh4ForEu5css5NGjJjBuQbIY1ALjMzYeN8IV0qgADA0a6n99h4U4I
60CaX9/6w/UA5TB+6q2IOIUEQ4cpTMlEB0NJUen+c7sFLmat55S5iqTxHA8DmH5dGMLNJyc9igkG
Jfj6CIxd7VWINoFyjK4k0RhFy7v8hr1EMcgAvhsVxolzdfVC07dYyp2UNqM3ZTt7rJHw3xgC2897
k4tZP9iy6xV7WgcDC1C4Q0KSklNEbqZIJF/Tl6Ce7Y1i/Gns8H64bsLbKnsEt4Dq49SaS6KARXlF
DMDSE2pHNRYV4B+YvgaVa5duzFuf2C1SUDKGSoNQqMq04Bu578MyesA6rH65IH6+TzNiv0oDOQWv
Mb8qc90cHaL29yhhI07m6avA3S7TqrAMgPLbbjEckCZDVJOA6VGSfEA/u2DnPAt5Vpvvp+idVaNt
KvyOm/W98LQoq1UPGGToTRlqNAELP/Boim3i0zovIoIBgrusvtPkWmKeMcSGZ4BDbMIinQRWhrjI
gS6u4A/u7GbNbqrRU+vY2qQCyH3OOkHq7hxSS7OQzLLsEHCt8pjmak2HrJtXgqkaJw+wRlsl/HAm
mL3frMKuvzp9Ff9tnZkYQfTMRIP5Rnbp0kf1yg+WVVJB+AOkZL4k067Hy42A3IWqaLeIrO88cUxI
P7E1N0yL25FvKrDfOhPlkjE+CI5aisg/AEUoczsdOs7UrHIkXYY/zGHB63j7aGklLygjsWmqCssb
02ByPumz0T5nm2WxQbCV/aM6OZ/xfINi5YFJftdNlplH4pnqUEgRNAeeovRr+isFbcA0ygvMtYqO
flo9frc6mP4SOuIQxbAPUET+VsiKfnBtsNaO7likeSRfPeBHIkfcS9sGg0uizBA68v1y8caBsX2T
xOst0GLoomxnURHn68P6G5OlXSEJzgMpSEz4oRqvRMibx/ULgakm08BLA6DDSVCsBRARD330EdJi
9hRgCqEFr8M4lavC0wsCnr11iBxil01WfBQQU8o2MXsruFKfvaRyb9RqZR4o0CcLOwDoDNqf0g+x
HNttUt6ERTfyJu37LwP92mMBi1bE12lQ7QlCVUFk3JeDmu6duhGSaIerOUPaPQczusX8j65dFXWz
ZmjGbqTjLZg/9x7iLAekthOJREtj4AsCiYUtvwGKZ10p1EB5QlAizEouywRVoEas9XI5Ayp1Pl+E
l+r4vMEl6Njfbh3A5NthzW2uw5ViRK5iZ5t43ouZjbLqTZQlsT/Q1TBlDQ+zN4O7cArsiWYceWyQ
+N2MkO80VRSsaCrQneaaJufJEdlUvc+VrQYkDKnvq15Hp7arYY3UYPrA2AdkqbyF0mYA6XXbGejF
aU8jZWEIUzSxOd1Yww86JRRRCIK+PcL1AalIRlOoCxwvpIwuYdnw7cuqx6mV5ojr74pxaKt3gMMb
JkdiuBWmB0t7UwMg9BANtD00HvdsP0plNrOD2XsLNFKAPU16ClFYA1n9li6nW9b+adAZVkBHfYsE
K+5BNz7AbVBmu3Fb7soKcU8oVeWAICALkL1mE4pnzes96UuzZmhTlChzCLsaXYq+yUtch+IoLnTe
SkowMEUAxE+k8OKifnc5mik5wH10Vs+QDI6w/Dy2HGs262XPrmsOpXeKS5NeSTXPSKLwhnsqOuk2
MatHc2/1j0JTmHSGDmpmQXLRnSv8dBDstjNFonJbR7oVIRD5yt+yU1UPmozivh+GUyz+RuV2isQv
s4gXfYpcEncynrXsxVH+l2BqXlyixo93+YOcEcwi04pBk12EIxXXNc+U4gszqWc7l3SUu12+T/19
qW4hH6Ak4qof5VYZDrrPwE+ExrdbiQzGXYvIkZhol/v5Hv6Enr6av2R8xckTnCBvO4gX7IDjKmDu
HkdiPsutzoC/mdMeEyVAjuC4kPs0hYptuKQj7H9J8L0JdVxpbxsmMiAXmPjdy2sSX9i6OYMM1Qjc
Kav4s1h1BFbhznTPl/troOvUHkCPL2kSVhDz8lFYm5yY8T4KhHW7VLAYax/xEkdZcT57vMzsMfsh
X/DA2ZxJ5qDaQhzd/fryftR2z6sQggy2Z1ARBCVEk8Fchvel4th5EnNIO0cvMX9etuUdwmtWfFSp
uaoafftpkWKdfUF9ryON/vJzrpRZpuOxbv5qENn0qrxOd5bzUnq6TEEHbvQGd/LR3yyOsM1aO23E
hOEvMzAtNHkHfmXxdm6SBj3VMXJbBBVWHfscwaqBu0svcmbT+zzxrnoY8tLrVXthgVMt3NF2ZPG1
/srJ7Iwpu6CwTSxyxblCMJOemn9a1iOwF5LoTXJWDTV2TDkjCdxEYgnz8SVY4imbhsVssLNi+pH7
Lt02OS1i6ao9ZePca6lVZxAjgKent8Eded5gwiB2vD3Muj1Nc40dXTLg27iMMRn4WkH0CwJ1OAJ+
v6kyNzsKvJYZS5BpWdrVRxfSg+FKxMroK943DYb2waWfeVAiehAAknkYP11pzGdt9TA3gTqj6pca
8/i2mYGmQ8OJqPbaPgrj5AO5ItEKfDRb6E5NjF2cIzVbZrQf0G4STfHhJboMNKfe5X3tRTwodYw5
F77aE/Plgajk9qhMWQoBroP16S3Tx3RzAL9cGzXZWynoqDGyljPnB5XgICUB9pJDhi4OUAxM5KJP
w14EyFBeUDTEPcUXJrQEFLK98eKQ+B9m2EVYvAaMaywM96AyTWQgZ5VWvwIHILoz8fCon2Q+uWLg
3EO4/K41pJGnBwIdje7bCm96X1HKvspccNYMgGVqqNOkS+WcAo67H7psGgpSnQhLiMtTfadm0Ml7
y+f5DebhkStycsYj8F16DAY2/ta0HgaUCMteC5aoNDq4JLEGMiHJ4xH9/dltW+PxbEK0nm1oVHPq
5BnCsrEp77/B3dAj4Y1/CSOoWcNTCnKR+Kr0dZndX+iTBXAJqfHVs6hQI3a4wpGGjWJotn66fDrD
VeHdg1iAfBSJ0pSt2A9XcTzFRlTNUulVDFuzZPwL6n2cCjr7PHVkN3U5xBly6MJ3wsXOegNhUk42
TF4mYwYY4DXGmOjWwbIPmprYtmdu6slYD3kUjfVcB6MIMqcqbU6SKKouf8S2AV8D8+/Jc/Q67MyX
sZ4QeCXpMlJ6mIMLJTNo4Y3yD1/VuniBlc03vdw1ha7OWeULZtXkN9OWxIpV8AvjJqF8jGl2eejm
NmZj+T2dnLFUZa/Of47Z2Z6oIycx4XtDlL+edWjbsebTeFyvU4yq8PMK9mbEj3pHjGHY0ex7y2J2
P620yi/GIVGOmr2YVTBdw6YN365E05aBsBSW27kUrJef0/vszqvsreSOiVs0wsPCY8lKVAvzNsFl
w9ilAadLvFV2G65uFykw2tmBb7Fm1Vo5so6fyjqYywwk43+AaJQguvj0uQt/wd8WMRsvyewdcsJK
XQ5rO57hy4wQHHcAuzv9xW7kmbPdIq5cU3ZYxvbwmHGrRDMdkea/J9tKE1j0TRigpFEVVk/9jDHA
Fk5X8GhEuaxda6AvJR79kvrT0GOgH1gq4Zu9NqkGWnQEtzqAIgEbLOHpC4IYVn6y4Q0H5XhiXWnj
QrZv9ekZRXrqN0VtTKl6H95nh2hBYsGq95PPSL6TFdwRCqKUxUWPyxo6RwBpafaO5/5NPbIO5Lvd
R4PJLfyy3DqFe8b6Vrmr9tkaWOvwbUlLrAu/kzPPe7Av4d63qa2MIM4vU4+VRGIXqWZpvLlHf3fH
cDCF//E/pLoN6yc768PM1Sf2Y+1xeLaRgWq5GWBc5kdSlehmUMNdryRhB/YmAd1MBWo4atkB1H9A
svN2qt7MNZB4Eb93jkXrTpGESsu24h/7/dwSdI4bEoLadvHJW0okAQRdOuUN4cUlxLx3XceqSyA/
f0Jbt+3TyHBHQBGpFwDYwvixMdlTmh5W70riDUKDTx2IL1+qFab7zE2KnlNiPGUWK+rgXXjlduKr
Opqk8w/WSzOE8DdX3JOHt2Yr2KocyFRQWRhTduQCA7cMAl9UiN1Ag5ddqzcfjH6eDEtwMQWR7rOX
KmI9jDG0nQVVOESd8M2n5K9jbhu73qVeokFJAfcmBp6vuFr6v7eGNphPqYSD77ZOo2dEKyja0Xjy
WL8FIpw1mdqpBeyY6qJ157ig+shEvJBp5bpswpw1ZPv7q4IJiJnffSfuRQvLs1PNBgEEfnr69UkR
PrTSLGCIi1CIthY1AG9sHSelLMQqlKKbZXPVrs/Z+CwEa+lB6KGlx6vwyhivrkWp6P7RRJQsFvED
VMtq9SGTelolHY5W31bREQI+UgI0owSYt9ygMRJXCGL85nFyVahdNZirOsO0/AQeDrlJfEAKttON
kdAZG1q9hfFJL1KI4UIfGzc9dMefOtwaRFNnKmNbsQHlmVO3Pxo9QU8RE+zVCXb70M7yGOPY/0dn
NtxtLY7eu68cRV0whGfRxdoleSUsHGdRdPgFDOvvWrw5bl3tx2OYqxQfcrp+vDgb5I2ORnMoNs7v
YEkUEzTZTGkM1MSaXGroAiw03rkiU16VIcCyh/svuy9P9AmrwuvBlDWdc/M7G4v7F7OKMCDDqjNt
TELV7KUD+FC5P+EzeuIbMzSlHCLAVh9mDw1nLQmcthqvcLZokB7dVJGoVXdLzhSFEJs20CTTaK6h
VJcvKEaSpR0YHdPsT4wnjQfzIbITRw1rI/XXUT6lfArfvLWE+b0iG+J+0LswdLVqx+LZtAiEvGLv
Q9WIecTNyBLgVqxcHh4CcroHfCTRjswBeBMKS3ucban1ieXHJUDsbEWFG6KnnL2Pe1xfzDoObdnQ
hFuBUtA3f3DcqAPaUswrAxkGFPLZgBTuBmBGIW/xHRs0FFDgllzs6Ltteqh0VWmnv7b8ZRsGfN8h
+nKlRtvM/6jQ7FeSuxbYruFnHgqnSACBDxosn4ck6STjVJ90PmhrNcbqQsenMcMtqkPvUhS8LwgZ
W3rhjLfD/0t4vlBmOLNXsJalUax7boyQKollDW+Dj3hYC+jbpJPsYdnxNuBnT9a3sVzYUrCTCZll
gpmMlkLz53KCgQ64OUA9o2MduGso3ZLCVOU2kdjJCAsnXz8wzIcxEQ664e7uRz9p9fjwdM9QBXYU
mhau3oKmc5RWyClIee4goS/UglAef+LYJyKNKXEygdjTVfl3qfBXK3VDuR14LPht9gvAVwQyDpfA
qiWzKoHyGPV49kjUswweVHVygkEseSS7DZ5TjTFaf2e/9G8lYs+KBW2fuRPXU/iD2yr0zZgthn0b
3XKJoNjtnp/SFWvUMKlcWV8GllYIYIpysU3fn3iGU4MaK7qx1n4rIQeqGQ/RQj0hpw/GNGjhLlVO
7MpXZmHCWwxENvelj4vPPmJBptnYVpMSp09LvtMCBhkI77XLUidUd76lBYU71Tj1ilrxqu61WE+v
k7/CxRFpt/8tW1DQrI+QO06W69AZHMfDUyI3CFD2BJFp3ZNb02apRz5FxJWUM/7Du0+8FA5by/Eh
SboMqmkl9LeNWGaSKNhdcKVt9hDRNzlDJ+fFlrME14XCZnJSEvNpVWtspShGUcir4M2ZccxJqSMc
qo5aVqaL9tRoRTixAg95afAfdMWh2BejwgTR4b/4dnEQ617ligyQXk+QuIBuwrTkHBY102tqs0yj
1+3HD2EOlAqcuwqpPWEGMyiN4E+gYNJPkqNHH4hQEEsrQYQUgScjDsXQlp+WyySdljXR4AHmKaJm
tr9z9Et3ecz/tWj3egd2OvZP5lH1a7g1k+VEuin2spa9MWwUGN1w06f2zm1mZnNOO4dZ8G/wCoqg
v+JKbrDB82l5lQmNgyjefPHDV0XAFVKhOrlk4Z6/BvsG+xFGtTGcY4YPvYUxoD5yagZW1ZfAFvNF
x8BfoMcbuLDXSSz1rnM1kSu2DfxZMCiOGtZryqzqjZ1UIJxJhF5PehEL+su5LdezwPVxAShBRLma
OIpM1e8RQiMDggPrEf9foo+HNzf9WuZCkPRuYYsm+8aD4bP9e2qQzNUEg/t8MZRUeu79kvi/cf/H
Gbkoqy3lKX6MhFUDoIl74p8E4OQi488iDTvCq7u76G+GkECOcLWXo/rNMBE9xB00VYkwMPxlY/jc
jGJychHvU+IYjvey0Vr+C+ChTnGFzpWgpnyF7hvA3rJ6u5EBxDIpD7oYsqktaWusPNSgmNjpHXjb
em3t3PrgUacw/84OhSiqoa8gPgFmEbjOgM6OdgmXxmBiSoKkcmbtcqX5Y6A3Gpz6Fw3h0p5PE+Ye
9NSJvG3dl5iEnod8prG9Wle1xthXywnfcrUM0wMNQrEiZjVEX0nAolN94pHYHjTA3C3PIEsvwxQv
qBVBjH4GinAZmW45LAl7qn9RD9pDkTlCqfHIkAuBwAvXVkveGFPoCB3eyNuTh0M/lvN1tZNaSA00
LLXKZ2uvIhizb1r0s8o0LlhRR3DqK/v2h62Sm52upiZlHLn/7/YgxQAtPKRWbL1ZzZF3YCseX+5M
9XgOUUJiM8NwcLk6pDTK6kKhFaYFHS6B9+q4cr07iaFpLC83MSWSAVMhulTwIlevCrYIjwgKeEgm
YTWVRGTFr/Tz4cD/OWr361kvpHfaW7LqU317YUshzFZtE88/nJPm2orPo4GXHZxMX8SPgz8eFY+L
2UcI3rXTZrZMtYypjQayP/hNGt3GOGig6VSl9GWx3iF6CRGcVNtWtgSeDkS4SM0ybBqQMvfuANJi
TgcIGTFhkcovvMQzOZkiLAJb4rkasy3E/vKONwzMFHKSWKJkoabl/0BHasa3NZ4BO4pQzfSReTJq
PVZQ/1BXWRSvMpcZhXF5/f8JFvWbbagTbMO2WsSnTbjXAcFfqzxzOgnMkoWJaivLH5P57hFNIVSv
MUioZf4+NSgcrAC53tofZw9auxUlHer5NMkJK9AS1lN1e890+w/RH5WyanoPhtdtWDoQxscJhQwf
zErujv7crmkQwuCJmSOsvMSzZWfBilEf+D9PdNu3sdZgUXIJyd35wEiPggT5Bb8vobxtte4tOH07
7DiMNXH/9xY0EKNfoGcEYORU7bVLDnLZYi4aznfFyvIDHuxBPOSRGqw1B1cq5X//HNbkHkmn8FHa
+GrRMf6acRh2ve5aqeMAfCbCTiUFrK5RYcEr6NxJ32yceOYrOcEr7wsBMwpDpDMgYwq36UlEBJgC
fvFm3ElGc17+BfImQQMJrCZLNeSUKF3tSrfxqGCG3XE40qgkhZb/m+ggd97gIn6zIAZhag7kTGlI
rralRtsOwsrQFjHOyBVXmF33U9CJQx1IQUhq09EYNw9MoohxFjrWgSpCalsV+DC+DH9ALAcBtnCJ
n/4WkMxSiOAR1hmH1VXEnlmd4IJffisaWrsgl9ijF/ZU/64LJlELpzLnzL2roy+q34NE/KzMtK7V
/BPaPHiGRW+iZJtQ0/COueJ/FlQSy+biDSt4VzUADZjwVZ20CwYgSd5hhlH++n3xhjCc/VfaXUKR
ppbu3p183Tqsvco9FYzX/JJqg1V2q3+4xSp6uaeEl3c7u7I7bSKoMBZz8kYOvJvFqSzvswRgVqv/
Wt+d5Sj/t0BPCQTvVFC1AKXwcFOVj7HEk4K3FfTBOlVnegOIeSBlWUA8/1GG+32k6iDg45dehrhb
2tez2HcarizNshFxq6zGZ6raB/FRUorw4dXFaOqRQM8sYJzWuiXxmcSSRAwexSnNc77p2FPsj6Qt
Yn8kAPdi8HfAzgoyxBjBjPVCRdYyHKbylT9LW6BYHNMYGsUOEGZiBhHmKQrJzNjM6v05PkLIPGNz
VNE8Czgf2Tos2jZQdyixBx+ZRVA2vCcqdbP8+z+K8R48GoC5IcPtKqyl4xw0GC2yMyEvCqEeH5Ql
WMWuHwbzBZ65flA8G73UR3vUCy7PJ7omi8Hgd7uLpkvcS+ptwRfC6ctxZ1aXX4YsqTG96NTUY0yq
Z8ncOjXnHPc9sxfLfhAeXSDqkAtjGxKeMxbxleesKxISbFvMEh7xnyiXVx0EM+AbI1vosQdhp3ug
m7viGQoD4NdB6x584d9cZJ/OoY7h1R1bBNdz3TUKvowdv32Drvbkt1kpSbJfRRIL6g8jYQAA9qLs
M0QFjJDmhLw3tPhVw045QvPBeKchnEhgH4KtFTj2MV6XoFZN0H5mQ+pu3DpaT6IC3igrYv3y6Zqh
g/RWVs4UsyW6zbpZSUKc2IqWBNdfWLJYTP/NhP/I1+A2hnI0FBDQCf22XYbpbKWoeptkyPdGQLZf
esUR4qLsqrb1W9X8U6uGSVOgbH0RlfWmzUc1p9Jt+74b9nhvKCq82ZpKGX7vuuM0erDPH146+5FL
dcnlEGXmI+x404sWYKzccIKh+CI1uaDloHixgXw+jdlmxB4AQdUTmaJMEJnC/tmXI/IOfFB856xs
TtEwoQ1LNlk46KZXuKbCtw058PrLGcVr8KoEN5CBep5SXxuZBNkG6eJyM6w/ErBCGPgsy4Is6IdQ
P4Sluniu3P0LqvJABGVMQa1i4dLiRkQazGGTmQL8rF4SJnyXGx5ra2Lh5oETABryBQN8sWjDlqwE
Y48Plogq8S6GxtufTE+882PDF2wqhHTMm5hp55KIRxBXfin7HRvHej8GegeUPW8X06DNSb5xNSb0
XGWY+fIRkIheWZmI/T2svBx3VA9dlsrQVObLWs4PfD+Tm7ogxKUR3pKEH5e5Tg0mo7zFD+3h192j
V0UTsGt75OdF392+bq7GWwoPo6JA8ve2CZEmoD32S0hy8i0VzKPSvJACabd1F2wFtntGkoFzaUim
eSoCvEt6VpBMaokg/c+TNvxjiJKV4Thq8sSq9Gb/osslKLfT2pNbQDnTSJAhL35EMkyxGiyPmVdI
z7da0GwBjeFlfaY5hOyhIfMk3BFTFBhG8ZEwr4HoIpJezLVLDoviD0QQIWZRYG4/1uq9SPnnWIEi
+R4hMgBDsSLiju9+tRwCF+I4fXUJp+7DGlRMd6qrvc4BVR0eDThMtkqXxdcMZzDIPNZADbTFSDNH
VrKwCevaYoG60J9Oi5udTcb/p91Cn5M5Zxu17MR7Csvl0oBqQ5MU507vcnziJQDYivxxgF7jwpn1
y5k78NBVDJJIlhacgBq0pFd74NcRsjxYPtVnS3BBlN/M6oke+0vhhZ6PTy1b92EBPHwGBLQuIZnk
gdac0Ye270gYt4pKLzIFN0hQvPsSZX9lXqnYLCqgS+jo+7BzH3LO53aMsHU9HaGFrm6JXSbTu4x7
zHry7cKRIJXLnR9ZRP8SXH9LU3MquxbJaGftIpiddBBPD1a9fatv31TkkmzRehoKBmOQg/Xsr2wh
/DRg1aP3yaAX3DAcJOoyEuUrabZTMAGQHEZqlruOCWsbZSJyTE47sbDXtlyaymlIXorpttz0A9ek
cfjvY89Pmx9xqxWNzWgLIlggfQCiY2zY6HJUErzal05mMAV6SOhsIoIIQ8xHqaZKzStCSOAtm/eO
h27sBa5u8SvzTPmiQzyDaGpzBNAHSmQ1wH6bEIxsqioaxDgTVf6wSzbZHu0ExNxka9WVXj8SP2jP
bsU+XDQjpG+C/eOkKnl42mcdZV+f/Z2Dfk85UBHVamCk9HQD0i683k7WifOpueuFgaoM8NvbUesX
wgrmilhuoM8UG0SX4+pCyQZB1JrKFxy9oBZwz/0vhQD1fZXjSr89rrNZZ3vuPIW1Xa8G+2pZRPwd
p39Vk4nvYJ5EBJ1XAYcyu61XGiFOAzxbzFbPpidWmHRUk/I9orLZPKhbBZ7q5szGCTofDiQC6Gfc
kvX1+CEOKUYoNVVf91h202FCh/lkjLnm1GXHaOrzaYqGWUcV5oeiww/h7PdSnFCEbnz94Xjc25Tb
HaN+20Mvy1SR5FyeqncPYX2D749WLGSDNrXV1g8bVBmHraXaCvWyQCcOIwWgqYSrbIY1sDJgac4H
Vk6iiNQrgzq5VSyhz5Ll4WC6ZD5NWxIQTxv900YUN/rGz0PkT/GxPpSZm7YiwXEF9tlyczfuWmPl
DIS/D7Pt8r+QdeTM2CzaT/Pqkl6rBSQO8jqQ0uR/7Wnp5/sMRivdu+DEs/QjUQHE/6yI9mIHYbi8
GxXcAZqyjDa3GcTI+h3v9xcdS7LkvF75qaw6cNK095xJpnKh4LOssykXLylJbkeRIuv9BpTIbNlz
8XgnibdS1kDgpactvXmsetB2suhweN3b0SiY3O0DrEbYCNd1G892/tjRj7CXA087WO3Xnju0k2iR
w6WMs2JyHwHlyTLvbhJRkL1GIpui7k6wBRNpmtUUUZyJYurbb41vxsum44wznvaxlK1z64GE5cTl
Yal5PD0tPsIrAuvPX4naXdzdVKx2XjFkxnQ9rTTTwwQB6cDshx+o/76aOrRRa1ZLWgegSplK/MIE
FZulvXIHtV/ldtrKXH45FHN5swgoWJAuj9JFgad0VvyscV2BNRl2xhxwUSbSnNDnKi1WPGKKiu2g
2ChQad6KPv/fpJ51ubXkRYmzF6LYhHalf8H1uoystngkENn7aIu9KVOIQuMBNRW6cZdBkraNhsa3
FNj1GzPv2ZCZHEWk2RH9yO9qToxF1kXRPLZwgn3kfh6WUJTrW+h/naax/lqXCPixsjy8R5ty9ubj
x4PRZjmHfT0nAQlYwnB1RifcplzljOEtadXpxGv+Nc4ttO0BnH0wdt3V5n7TlV1OxnQIJog8SLLj
eDORZwRlR+pHCRLgbVKGdEN26XhHmIzngB939jU7AsHtQunLmpEWpqDjkN6YTyWw2E0C52ljH6YV
A4CbNx/X5Sp5bNrNlCzu7+FsYbOK2ck7fZ0G7vfpYCtuRnSqo1+IZsg2/NuwzFxK4WZxEmIZRcQk
yHw5ybkbqC3bwEHJ4VOi7k76ag+IghkWp4Dw2QPKC3PXxsEIbuPs/KIZ3Tr7l/HYNg0Yvhiw0yXU
8ZXulokhxgeecZsSRWL+61vo35LcI5A/8TJDUUBZYAlMZDRzsdohQvkqMSGbDo4mqFUv3+bDY2Qs
Qrvfd0KwRs5pigAUefzM70oAGKmJKOIyuvnXo4IbKVGHU8G6QBVgTivQfElqSZcyvcLoigOlpZwf
V7kcE8Lua8/T8BDsYtYqnkrllaEAYdxoX0DRCs/pZxIOacIt4cZ7EZ269woJaXqQoctKFgbFNcJV
c3uA+2nu7Cj9RDDHE6fOHOyDSOSplHFgr3PzDPweplo4zdIP4tN8XqlgDBIUERGqP/bkcpMXvZq6
Fkjetocx7soGICvEBOlY07DIyWdv1oEePMGzeSOqVe6f1oEgUtCgYtMSXhRgssY1LxGvLN8+4Y77
KDzuSg/uv+2CPD+/YWqfgQoeEUFwF9mM+SvGY/UrhZqRCdmLyZpe6PGVwS57HqdmzCTY62WDAdjN
6eq2xYcUpHUlrnfZXil6SOmWGfh8nyng1I11g0F80vhb+nbPPEC+PkBzBuAmpzs+zbwV8YPJII+L
1oFX2Ohi8PCNMjdJ7FdwLhcgXny715GDAmV9tHsvS+rx3nVxnTDyqOXnNj2VZOhMz/oJV0H5zUIW
r0+Go+CZ4+pUpB0Dos73gnuOQwrCpFiF+VvFObUpdPKEmoDUac/yYweayMG3GiwdQK+LMZe4Y9mj
FX+HJkvaA5qOQrFVtZ/DrlU8KItbNwDhSh2zFZxaQAw3xg6V/uikrDrHSAU4MA7Fjo76EpMZe/qt
9nJZ8sBTZe8rSZ9Jo5hsCcEbG/lj9GiyHYgu67vi0D15WHuFe01iKxiYGXj6ZNvWjiSGa5kyEOmo
EGL8Osu4TGbLKw2zx+QN5K8UADVdbOl/f6twwse6ZLyi8p2iW43zPYTZAG7uAhfbBm8xvQkQlgfK
dBTbWkkIJXlQbmFpSadZqVYYLafRAPZk14POtYgx3SZagEjnMPMLLmv0HkWIR9By2UShh2MH3ZJX
LPlpdytXbIxIUtbrOiD69raaQ6g3VysPURXBkInfogZQi0dc2O4V5PqK+hjGaDW0Czx89QKiu7mn
kpw4VGoRWwlDb8rSN/CmlFN/Lzrjy81rYUhewhy0L6zhDO0CQdUcXTTX7FoAzKdgCWIHG+Lz5Q2R
9aW/oxJzUzWzzrdjJO95rKQx8Pa5DUyueN2hWtQVgOx+VmXJLX8GFnPP1dIYo2OnhczeqyltEAPw
9NCyS958RXCyOUqu+q6cxvIglLGCW5GHdz2eAqqE/DgSn08zsTaUPKFk0nvWONawztFLt5ecKGp7
cJ478fv8ebzEB8FSjhMorp3G4oSafgC7xWpbkJJAmKISMB16RXy5S0XP7YpusdnemLztHeHYJiI3
xak2lfhcxx9jddVPVLpII/ls6W5xl2X8nQcAA6mmQmgYLgk8LWRDUMK32Sl28xX5c/QhibJA5BSf
VpmLgHhGSyZUwNWeXnXahiqiCOpbSwQdnCFflZp3sNbE3RXTy+1vUxSsaZIk9O9N6WXZgztOBlgl
ejaJ9ITfw4Ov9EgsxKNdA/it7RBbSNM+IKcpfZIErt9IHRAa7O6oHS+JcGzPcK7C2AeLdJwsbo8p
x1zofqeCsKvS1GCvgbsXnfM0Glz133fyakcCT5jLSPlx5cKNh1eU6azI4KigsZ4hEphqKKjLcAy4
oRluSBSJpvJ0fGfeGh+hN57qbB9JANvbpXTQ1rHF8qMeQrD8N056m/KZOXnka5dJrEh4MOL1uHeT
JpnoRs3GgdSRnWwwpvS8HdhgI5+AOKjBOxR4OBE/JpBJuwmnZg9H3WKRS0PfYH/aWfOvOqP4+15Y
GApF9ryXi2QLmdnBrY7Ijo76dKpGaa+6syQLpH3tG+QXgEp1ddnbUvsVqApjfCFLdWgCLIp+0iQH
HDWyTm/zulOKFBvYD5iBN/3WEYb1tlUJ0gnLh8+MZZrJRJaSHpWCFG889jN4HkZVpz5VcMPv9Wpt
R+EVZFa7QJmr0gBWj0Kw61ebF1lNdjqwWKXGlVpBxs76S8SFCG/b3PXlJS4/AGb5SvlOsHeEilpa
+wh3oxCw6mSpF7ce3478svwAAx7v5os87WZHrgfauo6Hct7ewOs5q0h6Fkz9Z2IoMIl/JQQHni9y
bI5LviLKZHjzDmTAhNczEmTAMXgNprd2fTPud8Cj2AT+8zNlz7sKR0eR2o8WFaSGmzCdle/d2FrQ
eDCgcd86NSmVO20SzmWXXAzqQvI3L0Bb2KxFoNoM1soJc3Fggl9kO2mDGTtPozCXviuDT3hEdXiD
H0S5g3uHrzN+ZUGiQVIrV2/zL3jf1H43xfr8ssMMEnRn5GNSdC44nMg0mZiSLIMTH7qeIUGCDuYL
vtL2aQutbBsfMSxg9+qy0JcFiB25frCs+64UmfJ2MbLIROx3aeXDVHUduSuZHOPVFlGgCAs8mTyo
CKAXhldaIkJJ80KGi+UuP8sCdRHtOBbLIiDmhbCyeO1qr7jP4N6EF1rDTfJhhpFD+ifrEWqMIAAG
SvIoefudoUIjMbLAMcxJWcPcVXt1Z4VLPnc83lafBiifVU5PuEr12SWz9zZdubNFLA+OaD3dggla
qmdf8KGK/zdOSUepmC6ddc+JHXcq2VLVwrDg9aWs1/p6T+5M8v1skZo9WIMNYQ2PVP6XPeEYrwxB
7q6AgSOd7wyqtNXiOlDJwY9lpTRbr40CBXJvW+1ZaIsA6Rbuh8VGUH7dhVUSKpdxOR9j0roE+SF2
vFXnLtlZCAb2eBrtsIJ1bbzIWufG5iZfDW/Oc5LddsonopfAlVQ9FJFusu8Tw+mjzjEHC074fdPA
I1Bt1726cOH+XOXbr5isWqob3eEa+JaWnNlMyYipdeRrvV8vntVqsrbB4cNa0egPbFY+Z9wBjWAK
WtCwM+0cPZXrqzbTk1pdWgieVqIAPwGPBrPH8tMYdghHjmjHhnK1FQjL0FCfxZozkCNGEw8sG0sK
mTx0FmvqfQ0u3s/avvyHJvSWKMjJTl+2jIetnjHQu9fxElmfIvsPW6Y7TfvASkEeHzoQ30fWmzjv
/01xcofqGUrIsusqv9YocgmB+qasjvUTAYN7713XWAZGuPoTfRHc5fnlRR+Ymbfm6M+ammLfhbsC
BCRJbPGY82uF2M6GU6CaR7Q/r/k8/R65EA3Me4Tnat1oisvLglmyklRPSO27hzuN6xeRWXbuP4hT
bCXKeBPdl9zk+FFLhTSF6NZYbnMWUHkZvqQDiSMG36dlQ7HdEAKSHP4u/G4mjkxdp/MQJZbBRujq
qoj7CgdsXjyFhU2qHZ8uqK3pFXD1UopeIkbJAir4TSInVr7hVjoOVrGUooLySK55G8bM+ymkjM05
Q8Y0LobWQiKo4EB/j2lKgLkFpFLpvsrfONDFUHC7s5MioUcayzj36azJ/+S2xj8GVSdevG1OyQOM
J7CEHQMqw68PCdA8IkJPrrhl3Bri9wFSSkftxHFFy1NstTm/u1tPQyYnA67b35efh/fWjwA9dVdk
/DabN1h8QuoNOXYPCvas7lpEFKkehZuszDYhB/C7Xhbby1g7B0gMDMbsONkEQNTkqy3wN8P3V9Uv
cGy+KYXEjKr11Be0XTeSl5qqHxnjExPReP0vRIy9kyiOnjF8GMHQzudgdDXaFOdh0qxsqesevhlV
8PLMouycUoMvloSgd9xfWwsAkIHjAkVhJ4qy9v9F6MM5R8ORvD21QBnD5PsxJDcNn9xKshS5FL/G
lV9eydt8BRSSZKf4JcqgMvqYcz3Ekw6+DXVAxSLnmVDirATiKqeFEf72UawTMr7IbLrbmHhEjd9D
uSzraFdxHQvypu+zvgxHLllfjrgeS08SLnpd+iWFspp3wghDItH4c955w5226TwQH9d9ov4RX4C5
GmkmyMaiW8CwjxWhnS9o06KvIo6srYlfrJQP/awZcrHIp3uqXk9RjmorFlq0E9T9BD1xkDKWu3JR
blLuVJMQrZ/VhmuABzZCHVSPmpLsBtbLNPEhaHUz3rR1RKOR7AGHL3nEBbw/0aJfuh0SM8hjhe5O
yzBcTx1WSu5WMRfJWqELBlsGai0LMNnDj5JNvL3iwP06vQvM5JB/CceYg+eqv/yznz129XeEBsj0
xINlAhStADI7cY4uP0DwhuzjCYS604HkYphGWf3gc5giUWGHJ7HEtcnBUDTtuWJhOMUGpV3gfUzo
jhX/4mDgfusOb/qh6cAIN0hD3U2T1q1ZmNkODPYqIrLYdGnwqRni0/C6MXPLk+YPjddq2Y3g2pTt
Ol/sR2nWqkQkayHCxRDRkwYTjzX8aQSdHYY53mtS0zM9P9FIFEGGVZYbDFEGDuuyVRV++itDVmOY
qdPQyojq5SMuJf/7fj0qUneGVxQQsQFv1bcHBFiG5BzJfuVOVAtsYmcM9YEZC7LVENAouaLJVU1M
KN4UpNAxP2YjnAN4g5b1uuTH0YJAhylbQXDLF70BKzfvVS7lr38r2nmD2XPEusKPUuqeUeZYv/tx
DWjtgJvLx9QVz4KcqZXUnmJZaoFl04/J8hlZMXbNk3jOtWSZYLSFKOnzFVduoiujIqi8cDiCv65h
CtTOCbZeHu9blP31u2p6leNeHu5NVEuVToraSllIyueZewTJlEd/GjRMfsBT99et/2AsVN5gTjH1
ubyIg5QjUxmz1PtZYxJWj29jvhyoWhiwmfsuYbRc7UrPbFlI4o+f5hjL0AYTcqfV1d7LsWTRWmAw
+tfhb3eLaxzGkhfFzi7ALeWMnlo+fQWqDWq/Ll8BbaDidZI/oFbuuDO+ugBaUqSEj7Fx8ec5QrFs
mBWOIrx1M7J/c/RxaaTOA3WCQPwD7yTsjeJLXkBVsZAynFOTFhcsZFOLq/OS+Rw6+T8fPlngBq5X
k5oBugCEPgXD0YA1nUe4P29nO8V+Jgi48fhzK07sLqaztRUJR2E3MPNIXXX6cPSVDoWtbm8K7JDE
hUF5G3wETj/akeTGpQNo7zEBm/J0Y4FU5ww83T4TXaZRf6U3IpOCvKEI/yCWdfRNLtsS9TuLdtsR
fbcOvHgE80lwR52H7d/1Zhx8NGLj1ygk60iWyJTocImKc0jckdxKQUOPc+gODw75FPZfQr/mxAVu
R1frWEFZvbE6nhpPAuwDnq8c2xrsXULckYUffjfuuAX8OMEWeEq50umTujHk5mCDPZzJ6/IRtg1g
n/8UHQQWihyCbXbAM4Lh0qTHLgGWMrNTXqyipL/ZbNAsEDp67C80j/JdkcZW4OQolf2ehmz/tKma
wr5H9hPEO/El0spyUi70Sevgsdwc47wje+c1kqP+M/EdgzbKqq+sB5m1uP2IJLfwsxapw6VKuFoL
zt89miTHnEr4UgeBiq1iVxK/prAdHKYuERKYW0d43/Qu0uU6JdJroOM5EWL3wm8YGXJ2DlCYLkx/
REI8TPKb2n3MvVVyOX4Ly1+mCkt1ix0iCzywXUTIsKeaXLBuMZooGweAGFkBMFdHJDmi3zy6/++v
bX9rho08uCkDFW5BWc3OT8NiMbwcuyR+HYgG0MoWuN7e0P2RAo9waiPmJur/IGIs/muHSbrGg64A
Np9DvjLHNPHZy/QfkHM8VdA6pRmOVDGYdup9siehqiCBF6tsGdYVTyXgLz6XhB1tHZTYk3JQugyf
jtjJ0CvtGLIrKEoyNW8nOUJXDGVZRWPxH2mmCEyIV/kH0y1miCrWaWv1vOwJkLU/FG0mQSx1zyym
3LHBZQrwdqviVhpjMyV/gPSvluFj0wJG94O0VN6nUSj12SDpnj505J9yOanomfjqjAQFXMSD8IWl
QFnpA+mniw0htmH4kTVfe/KRvJho3nXc5ZvWX7ObuJk6UCsBW+gS/JV5tHk/qv/dXPpzvnslacMh
Uiug5yqim9DrxrZ0D6QgJTxCFOrfb3CmLLuBzBlk+5rofRAQeij9FIXasVioTjRBOTnsm06JC/QJ
c+VBwrqrHzMUphmqIJrJkbu6eze4Ll6oUWI/CtW5O66TU+Xo/hsg7mHTIXixDHtnen3ranJD/mBm
eDYwG4h4JghcKlJyep1UQJcxF4qNbzq8i3Sol+cqyzomu44S+dBk1eWinracx2HKqgjkoriDV1Zi
EcdUlSoBoV9zNNJvIhwjhtYHCmiGees0IMFtqNtKzwChr3w3ZDyv58qB98yrJ2FPeC0LA3GzWQ/D
Pe2PU15MTtIZHNNvu9GDBHH/PNFeDYNX8lukAZXHdNW4h/WmVp7ydF7+RfQXm3C9AyaI3DU9L28H
8QpjJobtuZvQTp+FBacDljw9rXARXnMxK/gmtvm5bv6Svi7IKMS9EETBN3SxwvbQBaLiJu5Ml2En
ex2+Ki+AgDWuo2RtLw4BrprYuuytph+zF5vvu92wGlvx7bY1vxws2YY+18b0XpCGoy72u3BLspya
Pj9JalpdsfMSnuPP1kVDodsuySZBAKCbhNhsXb+B8HY0gC77Ti39pYfbz60EpuQx0MQX6EtvlL/D
z2Mw8Ll1Y+AMkdKfLY4jj5/g6p8Q0ofQXPy9eHep9vpF+IVPxlOhr9K33IPAE7hE+AvC4U2FYmU3
jErfXUwMsvfeSoP7mzFEmPUN+u2UFzRqzqB34TEP9JKkuNwPyhCtXVB1O8i2QWPVzp53qlKiE1G7
+p3fEoDCdeeab4Rxmaty36Bb0NbDdtvQUzvGodXc+gH9cFdyScyg0YIpFz3K/GIxAlVbinPacQc+
+NIRrsbufiigEnEVUDEjNRmmV8qQbshJ3/S2L8OTFgEzK4GSiN8M7bxgJono1Bp9YQxB2qjiJB98
Azd9hAo7B+pVqOR6skeS9R07ORoV6JMZCqoTjLR2P5ggTMFyZ9D19OKR+MdRLB9vvqJAxoaNtx2M
fhQGlNh317p9EIIFvrPh4E+hGrNL5gy7qvKjwMcfU+WPtfwNzaLQWSqXXaQeM0WiTgJCgAPwMvyz
26Zwhol/Cs45ZcYMgVYRsLzGSU1az5WSl3+AHrjo1urWhrTXl5NuvV399ezXkm8BAV2dGLGHNml+
2kSl8T1xPGKrdwMNTSAN9QTtCx+lq2Sqou3Z/DKjZ9+eQE1hYa0qcXd2p3R9ig6t6MRShtNkZLgb
/ZhRYfw0LF/8y141K0mRg7579W9RJIvtKPoyn7oAnWGEjsGldAXwC4BiLPdRMvDmAZLvqvzOSoft
MkEdGKAFwz82ai/14QjRomJbZN+XDmfeYkQ1EXHGEojiLG4ELl87MLb4u30vOKHvVvLHiTiHEmom
XurzxiOD1IILCH3mdBCDqMleXMJaS0iD8cxOMmefAfw8/3RDOZHY+oEUByItDd/9Jhe4CvlJL9xe
cN4uSektzYvvj3rwFn05BUgTy3SkyoPZ0ncsjxsueGLC5rnsmsLh0MOurYQVfQ9AhfONEQrdSFA3
2TEDBGf6fl59G0JSI+d5rpt86mj84lxjOobMfd8z/Ty9o0rfY7gdVxY96G74a4p53dH+OQDeN/Ev
DRFkEOnQvUPuJ4Fj8LC8ww1zJnFIWs7D1HLDTVWD724qiWOd7hyIAuHUhITrNsbVIQcNCTAYKivz
+iIcbpUNllF2FTQW5UrgPnC9aEDWn02b5UC1xonwK4oriOKZMst8KeFc3pThyq7fu/mUWJ8q5/ZL
52MGRVZTtdIozGMmmXd0t9FLXY6mXOAvqOPRutWcJNz5sH4L3DQab1wwxhTN5QgYN1W5ZFjKlbHl
yjoOsC+QJlkW0iwyEljIp5P0tOWSO514wTliW93je8hzpPIOiUAB5VTzeLBW4A5Hv0737/LX31GC
R/hO2yk8v1K2ypTkYBb9PbI2+Xi2AWupA8Rya2v62GnLzceelJzltx025Zpdlvt9MDDNqRGD4wvp
BnEz/Axzplvm+pZY1KFSxzq20cy53i9z1Zfd8E1CDipOnd1K6N9lXWYyCIFJZIGR1FqoYC/Ifflq
H8vBasBwkEZucJSL1JpDJ53bU2Bfk43/WrWBKBVedTD1SJoiJQZta2NWEhTPdMCfAI/tIpLKrhxb
R8RblukPgNLvBY4CyOA/+ohsXtENzONpmftlNBb7jU3QVPWBAlpMNd0bhRsgNTzmCk/FAikzyXzT
m458ZSBswUlDB4pN7TpX/WgCFGmbL5jR97P1OcQc2iFDlR+Ms5j9FdfEr/rZSnhcZ1CY4kML3Hqr
cPv9sTRWomweEDtx1ZgdMUZotDNWvjXltzbJza1aNC25kjOOW67+b9h2XkFQ/3VAUlgVRHkNYQcv
2ioeYTb2AnUnSBODVjnk0AsiAPdy1teULgnIzPmVtkE3mdnsaMJwsHOPEkx3k+F5zf/cgOW6rY0b
DST/dx3vxKwQZtFNP9D9zNTZM4BeGyj6lejc5LyaXacxBmGvD+yABTL8aChw7rxtRztW7kDFDlK4
wlsFRtT6A0IF61k7maOw353ptMEA/VITNJvpmSWjtz9FZ97nRrP97xW7prJ6Bh04xySilY0LVAP0
uueeVGsWr22u3feHZ0jAps83h+jfIbiavjfBLQcLqMyFLhXicKfB9uraXAOIooc/Q09BerAquP2f
lrh3IZES5vKzmGWfKVkFETKj9P+8eC6MBloB9XK/ZlsgBKXZuzbkb0XHi5Q2fD4Epy5zUUJhQZ3f
z1wtWBIKdpM9LlBl9k2mHECnacdpbB4eybFWiqiLgIscU+UVYXq97O9p14wsBjJ39eLv9s4+aFfk
e/um9IIi0MAeId1V8M+Kdj3FEscNRV5rYEU14Gm2YQ0sRtTzdLuQwTrSFDYAy7njYhaziAf5C4vK
OEY6YUqBU6/xsIxK6PVr7Q+RQtVJgjfog6gNsfOOA8mAEqBOvzBgBcQjz0Qgmh4jbtXg3i+iH+XG
Y3PieUrod6kmJ9Hb9zuMrA0HBaJoNeh8uMWBCuJSsBtEiWBcu9+0Bwg6piMx1lIS0qDdSTV/KQ6f
eFIF03cZcNe7aE20wHh+bSfliMhheaS76qg5/s6T9W8NaOIT8cYgP/4bUfhJw82Do5s43CV6aCpH
MfqrM/DQwg3aBBG3wKvxZS29Yh30LOdvBEBgzhIsaiEWkrWC4KEJq7FZcuzxlsiq4ApoOsp3ApzH
H2fHBxx3vZE142y5cY74rQ7//hf9FK/9zv3XZoj5lUr29cJWencYyktT+tugDojeVpPKgT7EB0FF
fJ9noAK13ggpHSTHe/BAXg5o/A/SDVUOAil+hbJCIdXc+HTAuNeanuoQmtXU0FdUCLmNVes+EGgj
Ggthb8zX3qC4wnyvyUphSzcA4jKYC6adAvZA4BWUFRzCbVA1t15Ud60IDK9tw3XYWU9bVX9ymd64
o2j0/0uP6V711IpxguwxY05oJpb1Rr1XhJs4dT+hy/B5oFwdjrUkEZ1wuXM5vV0dkSZUVMF4v7Tr
Gq3ZktnWLVpi0GERDeeMbALFJqd2dYPVuQDwvB31nZhIsZDahVOuCPxq81UySJcGZHOC85dcY4Q6
8u8/y7RMw25JJN2z71I6h4ed9VDiBapc1TZOV1I6/ThzHSlYOUDF60Y/KT0UzSczJggbX4yFRUgB
1HvAopWd/bGrXU1haphaADwAmbCQpBtV5YJG93rikvuWXQ/ugApwu7ExsS/YsHxN8lHQuJA2Ofwl
bPuwNxePcqoEsaozKu62q7j0uJWBx7mYOAnteYmq/URAt7rBMZaqW7WZwYVOcr/q8GvuvzJdCAvF
ai/jVpHCMOYdUUqWecULphRHJ4YGJPBWPg5G4SogZdDSpHAr3ap50V6874v+0kBZkzu/PP9eabch
rfb/fGxp4JuNNWNbFSiMGlXqyowxItOMGkAHZlJOTl/nPilnS0vMkThSIDYKyl3pcGmofwWNeNMl
xx8/xab3Kf3dfybP2v119Oz421/AqJcLONoJJnggGL61dAk3/JCntKdd3WA2onbPBnQR2bV3rewg
65BL0MJhUUBLvZyiG1YlMSAyyl7cCCnCcdixDml7nbiJQN4PNbq38+oVkOc9jqpT5GuQU1jiFDI9
DWkDI2IDt/H2sAsOrSiAyti3biIgl82F09uDaOPLmhkEy79HdCd1qrJVMO/XM5e/x6A7oUD45FxF
GCk7b0Q09/Gyy8paDv1uhbTgxFfbYanOJJGAVM/nqi5uvA+TrskKQxvzwzp6EQdUJ2+zj1kKi1rJ
9+hkLPZNM+cUAa7HZFDHqZV3nDo2xtIrptIOxhb+4ONSQ2UFXSO5TI1/ftJTN40t3M8BCQlLob/z
kMhMBdM5IiXDEiCRDpvTl3gOAwjHZUyqrLqT7QmDllqJ4IqDgKRKRCxJZSDMQm2mt+cslybFM/Y8
XOTtii1EHqRUYAlRZ+Pxxn4ddP5Y7kcZ47lkR+HOz0T21t/hvjbVwgnjIORHC5fw+JrTP2GVgGMF
ko27S8FEKjJyVVZbVcEC3yC9D45DMp1X4075ctORalYIfOh+9HNzgcTbdugYmnxMF/4lQI/zpJq9
MRyDdLs9sn0Kb1EE0eoUD+NlpAh6Q1UA98Dvw7kT9nc1d3qALPeC3vC5nL1sAlHakhGNJrXXB4k6
K+Jgz0SAcJkXnDS+uAWlClpMW1gbXzRT9zpioOGs4FDypB9Z4ivaM1SquCS9QAS3GcH4az4Pw7XN
eblsegdPRB75HYer188eR81847mazCfOvq/uhAmSt9NCqU526wYO4Pv/ksp7s3eya1NWsUqmKyxB
RuYSD/glNf+C3GoY/anXv7WYyTdWeMnMOVh+TExG9OJJ6p29ELSIzFGahf0hNTSIdPc0m6p9O1q2
2C+hJY8OGc05CDKBzQcfFqDcIpLi1NQj3kIbi5fPjrTa3ET2mrZDsCqIkudLaWmGRVNrPUDmgYMD
+hDoduhO/iy8IVUfEKnKcRRGbGWu545acWhCHivAarTJgde2oKan4yfkDb28G/BLBem6/aKSMvzt
YiExpMd49CbnqiYkQSFuN18/hKKKhJI4FUorJdAywiJHGh21xMKx17T9FWIoRu179Enua8wYpsKD
dedIDyZh4JaoTUHPde4DrghcilFxq1QXwLLoRneOJMBNwdwTGQ2PdQc8NOzksrORy++TrlHxZn1A
W9NWNqxJm9IDTAhO/kBc04ALDK2H6+VjVsU2L9D0PlsQPjr2CzmMYvO69/NH7YRND1qRJWTonI06
8JM/BDXfT999Eu4dvoZTMLFNKJid6gRKuAjylVMEs4CYOv5fm+fK6/iMy6jOUac3X2POk5rn4Bf3
tgMKzSCE4nncGoS4z+G+Vxf0FblV9w+RgJnb7HFwQapEABoKlt23uijjxj2Y60SFCZJW28O/ZGC/
rHwcAo7kWgsy4ipp5wxGhFa9M3SxpaBZVZ9EdIUlEWD75oN84RRYgrMCYuZbvc4vaMjkb134to2P
ivPZQ7/Z0+UPcGJle2DCy8wzQRFJi+WFcuXa/rKhUkl7XgSX9RX0mjy63LqnJNp6vTj6ihRJZQKl
I8GjOEIAmBnoq6X7GQcWUf5b/x/kW1VCNZq+0mdZHlgBF7bawCRaHONXaIFDzP97ukC+wdueMcCX
C5EiGhtPad2ETLj7mv5u57SnxSb469vGHh2etwWUC9Roi8P8K0pJtEwEjYpH0MH1ZR+KdGhH8Ne+
i8gWZi1UCA4fkqN2YnXNc1A1kvgU5tpgXEvAqjUu7bY5GCdKhoyrKktJYJZSqILyyazMCrt2IiiO
JfA4T+O9Cyuy1MohSd5XShHU+hUGfmZB4kfE+7TcosGJ468d3CbfC18CoTqRBYw0gX19OGfVU+aI
36YkqAnbs4gXV7SouqbEqKDgQ03KALyzDiLgHFhAzgygLsEKc3LdieD3IbjN+Eb+PJRqGPCWBDk7
grcSRJa3Z4h+PE524LfVIoWsjGjKiHYGKqCfm8nBoVqfE1ID6Gyg9okPb1QMV5X4zDzLWm7JCcZx
7Hqw3uxuY/oZVJNWMCePNJ4gtZ3kSN2x3zorVFOsEE4D3EFLLBpI6zwztdWWNy66WA59E+b8C0KO
JeT0TJ6FG0UrsacEb9AfEM8PleOpsm1J9XDaTLXBRfnLGDEo6i0YXksIURLB6QfZTW2+1V+qcWtS
nqP8noCFUC0v5MT65CM4+XQYSGM77n7hD5tsvLX1z85x2CEzdV6GLyYglkv5MSjTZFTQukxHCYkD
X2iK7x3o0BFhEYaLCRfQrOOv6IIkm1fhoY+sg+mEJqoEYgaitH7wtib5fJz5T6Pg31xuvHH/7JwR
Anlkbzxy3aSpRea4c9jvwDzL2Tuq1/wTS6AMDDUtfQMAEMh4LFoDtr9wp/rKRqbI0zgdysctS6pg
bzDGWFJ+6wtgDwjNxwCoTZdsqsCJmV/JTLW8DZOGXkHXq+ov1Fhorz/D2Gc/VjlTbNqKlEVSKvBu
iwnbX6kZ/QoBdASro4XdNQ7vSldhLrVyUgy9AlyeXnOzSyq9u6LTtfccVGsyxrBu/dLR1FwRr7tB
cdzB5Tgjwzn1zwoXss64F1nu7jmIPeSyvqH0Gia+dTMExH0z4mzCbOktjcKDqj+CfM83sOZlnhnD
1YMZ6GU046rr78zcbK4zVRG0kYMm/Zse1kT4zpylOgZ07hvL7EaZEjWbp4dH7Pexq983ddqAj+o3
XVg7pGIFGdTtbAunLYQ2yzcrSEftZouLRgGRm7IhapC4+BA6D12LjxodVi1x3AGI0xpIwD2vPQB2
ZYlqtoRr8Cu2frvUGR6CZBo62f5daGRIildI443+8FFDnQVTO4g9yVol7kEfYWabiL9J6p9R66BE
4eZMswDr24Rkg64QicOeHtmLsLTrj+PXmz9brtFZiqpvA80qed7NyVHKY6wPSNkRWxmVOjSeNMe1
ZwUXGVjpfFvIkps8WeKxg8I2pu/551WFkw2tr0Ly9Kk0eN1xBOnlxp//+emBZAfvygSwTX9SwbUH
1Sy9XAi1H/WXm3+daXZVkp0iaYwoa2SJL06cTOK5hiIs3wQ1ZocQXixBi88Pp2HKHl8iCxWswqVw
g2luBE8uTlqx97c3Kr747zhj+9Kj3Opl8r3p0NdMy++8TA62mMIhOstW/hayd9JWvu9/DCDNYwO3
payUUXsE8B1mp6GOuBuGPkVxKuxIL3iSUSDy60MY22r9JK6eRNe9TOu0yi4Aa4RGn2D5mtJv0iKb
/EJt+hC8JNOlLcSFr37azrYHWQDjXSuVpZL7Eax7RyzTnammfdvOlFkRLmBZD5joUxuRMH74cPVW
3ay6a5+GZka6TQ8gSobw/ccFWU4Uv9ohkBP9yKJ55QDQKczQeiTE70L6X7PNTQ+SFiNBMU/9ZS83
6XW/QtuYLiOuNlBoGJzjEi5e4mUx+T0wf7FJY5Pgc+6VnnFLzVHYGkRxVmdmlAZB0GSbgd0Di81B
p1uw6ZCrpTZw9fM0IiuEdqxRbgvasAf9UG+gbUNMgwTEwwWACukzHxjWdxyJ/kZi/A3Q9/MNjXom
sWcvEojEUw7yM9YeQ5Iu2sNbtu8b8YLjcR2tQ7GZeZM+rOdVf5OT/l9MkKSeOnEP4YMgyUhRbOUn
2cTipsDHLWn/+mTr9kYYsiCjL8zfugtxis0tN/QZWq17TiGUQGaw9LKAP/nJoeSsCePHWq79lhKM
1ubgHdVWK4RtsGUg/2MJ60rXoB529JEj6tylJjD+HLZ72UQT0eYD7eqUFWoBLadTZCqYYiHPRti4
N1PpqBgQ7bJp9jnyapGUVvtCojjNeNbrejYD3bvt+f0qUq2zh9GhUIlwxmEYMIJ6OxjPK1mv2Bqb
gB57ByO+gRpJHG8l+4OFowrwOa/MjUkJkX8GpPtTl77MHvv/WONptMZQE0DIk5ZXMEo8VAa2AY/p
51xmWgAxa8evgffW3wueNe48+2t3/FAP9kZHY3O5cl6M47m3wiHiGZ2Mglq0/yo5xKbKCsGGZ5yc
iG40Iz31KeKnUNK32+tY0bwkGcBe7FW/oPVsyCiCgB2X0K6tNgC0OwD1Pygz1UeS52k+5vf8GTYA
2zY9q7SvT2w259Vble11IQL2Az0Pq2k23OtNnZvXnv3zw33l3/RILlxel17PyyfIFj7EeOPcLOTo
/3XjGinoSNxsgeVVJgJm+jtABjhEQlf+WIG8K2sljMl1s8/EsDgWX0H8HjDcS7+jQEEtXKeS+UZm
VP0xHCGZAdB0Le3MjGxfmo5eCRU5WmxOggMyFhamvy7QFNQUddkT7VPkh84J1WYJKU3nCgmpiIn9
fonwSI275B/6Y12jEMEdaJLAzJK09ZMjunZLsbuxQa5/GCJtO77UH2FT/WtU8y5WVOodw3n1MPV+
NO5ElFnE9e9dai+YgPeYOSQAChG9vRpU4sMOfRDdXDjvHQ67lwr92o73lPe0ZBFnZ6CFnus6YxA+
iVaErukMduFNRKEqvt3LwTwpHfazcjPNCNIJcdtQwUGG4FYxLdmIffDyKHIomst9HlfM8qX56Sai
ptj1PMhnLluru7WPafy8jWA0BpPpxaA5yAjsHaeMr51VTPQKwY2aspBOQ2nCv+yW7+x3e8fKeNqY
jWCBQtfL1YKi8n6Ri6aF/BlShcpjYuAr2nE/ogMTNXlyOBngDsTlalehsOFObMG08zj6+5o1xTC3
oH7VW57yWktmNEqBvynh3PM5VEqWlTgzwQKxPuuwAvx+NeB1HC5q8DKJr8XJNDNZju8uoql4J8ff
PTqXYGy7hiR/Q4ffjOWXbvpXiGZer0zgU76UGoH6E2K6hEWIZt8c+Q/Ly3+YfFd2meHApfZMWwdH
svL6wsbHzGVkvWERFqm3FloFLOsQizNcH163J2Sp9peP7wVYaAYuDVY/6Y3LkmlgzK0NLuhIzA38
A+9jR/3Hwnb82VR7pcFXj6IzW2/snMB4zwZmUSjW/vIWZqVX63IkHCygR9UynK1MWE4nrWyZLsV/
8LLxXGfxMVfY5GTR6+VIKm2GZIwxijy/vOv3SdwjK7uyYw/ltDSJWlCZFFrzgj15b4yMu/+uGMOG
xKlDv9CqB9pOQO7w8q9cNOoD0bwlzcOoz9LYqyLt6ikfZ0tUF/OuCcTxh8g0qhnNG8vz8hm4DuiH
ltgywe4Ht9zzcFxsr7CSMQvLTIOKJNJehF408foRnLO0Y0tajIOQ+TJKlOHhAtkORT1NZnQ5t/I6
dsxzg/Cd4pLw1amFjQZVMD1oOgOgbW9pIrCyGBeBrYAVIIY+/P1qouwYomby1YhgXFwA8/R5EZpE
IOcFqVQyUZBtZQHPj5VwpuAMuXUwBqMDCYcrfgnSwn1t8eD8oDJZ1MsJ9mUvFbTWJmdVWaZEYqRi
0IlG/QQFW1QBv6Vdzj6v+PITfesKanmXbU68ydNm4WWwx1zfdrm0yzlyWiOPAMzNFCzijhiaazWT
G1FnXHLUc1BpXe63uTEVO6xZCxKrZ0/MRtWDuqLCSGt+OKQBZE4P5QaE2sVMdyJo1WBBgVenmD+F
zk9gLn4XYh/A5sz1fV1lQ/2y4kUsYSSJmXpYuCoIfuKTPsX/w7ZxbTu8sjfSxvmkMvQsCWGj0t8M
mkGXNy3y/Jbab0M/wWXlGp8QZKv4Af5fkbDF6wmAUGlDvAali4S8gGh/ZaV70ue8TXlJae3OjYZW
jRGsvi+UU8J+eGZ4TlGk85wjjsoxcV0rXnJ2bh6T75AAUu1zo41y9jPqXwolTR7veNJxK7kb3sXi
ny22kjAnJ7IFQuPKGFugyfoYofSHG8tlXqy6kuo0gtRfukSx8nOaffHvuC2U0JrFYCHQ/D02Hxg/
NAmovenrJKYHvLSkZ+f/YdZj0l02+7sHLsH++EoAoFkNm5pkJ9r+CA/6vXJvL9retfFdJgziSfyX
JC+I4vJPMNwTvsQCcIN+MJowR9gwLmopSBPAxu8RrCBEh/yl1HaKOzKNaaVa8UKvjJMLdwHIEBrX
V8FsY49Os0/o+3Nuv2cO1V48x09XxdjbZD376s1cXv75Q4+y8N0GZeudtzbGFm6ENheFmESNtb6m
w/3ENJXzWM+QcGMG+vPf6BIu8zmo5/Gbl+1kb421rAB62olUe68G3Uri6hrjsEXAqF1Nw9ixnb9X
hJayPMg0GO4i7nojldt36XiLuoOAUuB7ZQIIyRFHd21Zj6cC4NJoDDpci+yk1jAbN6XOE7rDGWu4
SocexlQTg8/RuxZlJ2ksJKCL39XB1a0ClQISGa0e/w+YJfclBkc6vgU2iKyWrKmXmadq6LTQT274
CIhgpeXAspet2pOMl6a8MFKZWiYodXh3huixBsdnsFsfbNev9j/Bk+WkRkNy4NAJlLEwSpgLxOSk
qyV5toHtMiRNMSHhsOFJE/DsPqR/O/ppLkIK+uF2s1P7iX72G0T6j7unwR4fn/MDg3Jvvzb+hG3/
RX5uD1MRtdrHibpZvX1YRDh/utBxw3f+sWEfYMYXdWN5eeKEMWvmCp5QePkvzu5aMMD4pJ/8h3Tg
7NJQQ8XV85UBDMzQLx7WLtdmJzUxQaWWUZqKaZFMSdbxRqvm9xLXI7mD/DqZV3gmptEbtzWLZ1si
rc+/t25ClLqW44Ayafi8CAjoQJpP8Y9pQwOHT0DPRj2b8gT+pnFrB/Lq0TFKaWg/Z8E5NrleYXxQ
5+wsatGVqchXd6pHb+PmDvFUojrmC48IfD5pSbw6ZTUniXXPf572PfOVuAAlkJtkoFH5TSDubLIO
GbBogvT3wqXTIN6WXhXPayQToUkmRxQ5UsKO7P3fnNY9Wf5KREnj/sQtDQeNp+wtzNY+PMY9vHTk
rIG3SJjokRdJ9wBSUE0/vsin/eKBDdouQpx0VAYkujW6A7ckpSiyaDr9aU5LccPExCBDMeGWV8kW
Id4VVL1ujtGofsddLl/i3jynHQydR2fUQ0FfmfkKmrpfjz47tRm8zDDCf8kR1ciig5+xS5Z7Wkvh
phMnJrdTUA2dWcwq/Fv3CR9iw+tyZR7ifqbGiBifsKde4hXU0DwZCoxJGciBm8j0T8Oi7fbosIfX
qmc01Qn7tTmak27PvvG+qXMos7gNdiBP/KfPm5cnfXwyupt7Jr6QBVGZff6lz3r1YqX5eDxmIZGX
/+r5qmxKY5WlvtkZHhb1KpkeAQ8+7zGkXdfajjNZNEwfRXVMuYYWN+kKWKtKul/FHiD/vr90x8ia
tWmRmjKkqD+zb6b3ipLy45/IJCIvHZew3dtmz73KRWC/yGOhltqj3KILLdwewwJgHz22DiSf1s/f
1UsBVZ72EPTlMITHAFCqeCTYmsVxja4AXgO/NQ0ikeBWhtplwNcPMKYM0vxjl9Ielo5VEV18vdVn
6TRwVAtrKoHcNl4T7XxmL0P201lGcB6sANSwM0VS3vP48XTyYDenc413r5eRAI9UBQUdGZs4mgdD
8uwrC9DS4ATY32eCP2hOoGKvPMRLeClYy9DQfReQecP07nF3pnvXVqNonIl33+VfWliQ/DvI3TLJ
jcXEtEErlwshYpImftp6ncU1nj/JLy9gLbRD0wHxACx6LvGoZjGzMCwrTakVd6o158ZilrwIql7M
E3Ih/BmXThTTLreD57jYRg/OaAHvsJheUy4BYIT9vS1bbROGdxoflfnVa4feyRYHtfqkZ5+Sie8d
bGd9hlwaFx5AejTSmTJRN0jqrKy2CjMcq4WTSIQH8Taui45m35f7+GBhYKaIEp3pnNNIp7nQQ/qA
/15O95sh5TXOqF+6Z8tlCnAChn9X+WSoaJrECbCpZDDPvqZKEgoW3fFiRfHwD82wfr79zSmWelSb
Qx70SNPhwlCaufz4JwxoF8k7qat5x2Mme1ffL9yl6YWxkXmDqL3K4SuN745zAu8XgVdGc9agoes7
1OiTDo1mFdoud7T4VcCyO1mwH834NQUUmkFuwmiAoTTEPHjWDV3YaIp/wXDrEVjdw99+t9SNYO1h
WKVyL6Uuz4Q0jP1lYu16ScW/+jb61Uyq/TK2Pkc5ZKpMoQYtFJbvFHeNoHsJ+c6wUeXTK49piZvN
rFzgS8OIumGTRPnIE3AjATOHeha4sSPp/m4db6lPPk7OIUg145naBh31h5WXjWkhYlatIU765wGi
DA/i201m+BZvHhmzJ04HuaTiQcZvspyNqlF5YPpP1AxcGmt6YYtN1Bh8nH7yFL3d5MQpUpO8l8AO
YXMa7oWc/UL9SF7W3BHO3HSwMVQhA+GVQ4pxKf2inXIUAxSnb0lpDXFGVc9o2hgvAzImmJI64dcA
7dZEpMvoMugY50FHjOvT+1sYbV8mi262Uthv1f78i3I9CFWRXn8xOuHuyEGLn0+0RsU9BdfVAitN
WvMP2W71rIbRk6wHEnuJEPVygom3nu52ZF2TMOeMFa8skFVn0uPZRefyJmD8zea/Ba69Es4gIiCX
LaUR/kIerY69CKCGjRaMLQ3D2GMqWXh15jwFWdFZy3Vn70110aqZTmwYHwyVxJWOqAOV8CgX6Xnn
Ddu8yY4ymAqKKr+UrhmZsO0+3+8VcAgcWvDr2gjHQcMN1DXXTnJU3S+TRrMMy/lNvni0pbz0jVAj
SpzA2lXb2iyrDi56/wuGD+uZ3Z5MO61nm9pDiQCm3Ixk5I3qb1PwwBk+KJ+AXszg9lNYI05JPqY8
HkdDoHlwdYw+7Ydd3NOOlZ4v5yEdpqKigtxOaFQHJxTLgW9ZMOq8C+vCz2Wn5oQGgkQhoEh0e0/F
E4lpI/SCAXg5mFQFfkX+QLq3rG97oAXCQChFv5uq+TV+8CCbqn3P2s2zznsCqSnvwBKClDfhmZuM
QdsFNLaSy140f11rFh8XqlMG6PZ6CEjOMXI11zO9SHYP6rFppicXd02atilWuJaxHpHBcleMWN7T
liQKXCVjXIHeYjnQMUZDBmp7WAMv3OxtjLEg6opg3WLEb3vqMS3xUcRPk/n3foj+hV+Osb30FWTX
z+lRnOh7ELN2prtVXG7kgC8kMcdDP6HU6BcCt1eWrynJK6KXkXIs/616NGJb3iuencKfzWHpuTxC
1Ru5ghV1MTE7N6PGHT/eJDYYNqY49Pmx3+WhEihfs5HOqQTS63KB8kUGcoIntiieMXtgDKqi49Lu
Mn09ABJSCSE67+R7pxlK4qr0hMbI/SwYoCyakMyoDDJgs0TqidCggvZlQLNsPYzBKf9Tbxdct6pb
gi8MWPOLqf9nKuJV8fwflzAHhMHupPcbAQYmw/kP7jEPDN+o28O0F7eFiufYw24SpRp3wfeKU3Vu
fcSRnjw0zAxMWrzOEtzOB6zQfziUq6lW8Kj+4kF8kCa30ebEzNjxtRT6rgrZxkYe3MVETwcMuH9v
QLKf/J3Akwi1xJ96q/aqyiB/XxiRbN8GuVs0ead0OK6lXE2WdqZeyRosRChtZA9LvOsPlEj4pPJ/
tkCFHjfjaWii1e2L8htT62KTF0vakEWgIdQz+2H+ZG1QzbN1s3bcm4IVpwg/ZYkfK1lYpgdVY+Ft
bNPUt6hAMbLczewAeIvsslKL7xU0CXhIcDgaxQEpD0h4D27e5O7vbTZwBWTGQChfgmerB7Kch+ju
Vj9UeI3KXrIMcZvgamyg5Kzreep5M+fPz2abRBLxMY7/WFSjmFIMwFX5KcTuZrrT+8hsQvtTzDFB
gXj9+HDojViM1Owf9A89pG2dKAqtxUHATE/kJVaEzStPEOkGOy7eAuf41Qni68R2Qyto2sz2Sk2h
HANo8e8piIoTK01JraTUDnzkzmllYNWkyg/1RP0eocoJVw7abxpESFBX5V2tO3i/3Do/BO0nqP0z
GPlb4VQBUBRBv7lt9aZEkfarhF2O3k+/zNOMO3UxurWKY7W3uNc6wFEWzFPq8rnvSaoWR5lKHiCF
UsG8+Ozo8rVi6q2X4bYegMKWGTSaaJkc/AON/t081RebZsx9CGao3nsmiMCe3gzgmtZhfgce51fy
KWm9pVGfTBZWDhWexWbXWwFKHsbtirOUd65wksYjhYatPlqJPd1i+uG8yXAsUqkFGl04UcPa5b/h
j16c/fOEhnZSqKm/ewLyJHfgqTye0HYV85tBbkkCNIy8rh3ST7PTUivI/u0yiTivBgzOR6/54tev
yJ1vIBgOvU237BGsgLXsCmXfTqWcIrPLLMWLX7iYCAMU3u3jU4B+MbE4xe7zhyhHd5ylEsdlqUjW
/uv60+fvcMczCjZd0aGSv26bZ/thv3qj6dRlj+Sdd0DfJsAmCJfVdPV10ro7CC48cYt76uwOZR3b
37B7sJ5vRJYevYwLFEsCQwOSPndwYcTGLT5uvdOrvG8wvbWDsk/41blOE/iLsBp9Lqfz0sOsTetA
HIKQwt0lbsu2+cP1OJDiOQzlwIqwm3ZmFunRVaYFLoj3UFqJi0//T1k33vGpHbcQbOg2NzvuemIu
1PCtCCLhTWmfJYO3fIdVETfWhtgNZEzoDSRy8qSrBqrvHPrctWjPWUolMfGt68fdrlDsqWdU5l/k
lR6ljpAV4HQdSQ854lXpxqdtO9GG+qXj+09Evytr9cmHkjm9PcyscB8pjhhabn6laZ1W1HQQXDKk
wi6IdM5p+PtM7hcsAxRD0W3sHwl0bB5p9fc+aBNR/B5f1KXcNp0JAIcMWCpNmGhB7N5sv1YvMtdX
AbUP95lI1kGVIHukPA79SuHrNf188sYN8Rpwgs9sqlkZu0SxY8Uj7uVVf4e6E6r4hedkukK9u07Q
zUvLlkXwucuQdZ4jGe523palqhT6SepdkDT2IhhaS/GHNDNldPdgUZnsE3x0ZpXfdSVbplAxSHfG
gWESPtK1q3owfI81ctncYzcHG+9KfKz5yLAxLkTGEeGe12UIZrX7V6CjmsoP6g0Bbtbqj5UM1zO7
TpYcWdpJ2gltN7aUY11xo2TI5BuB0R/YSXA1OlmZMzZp250WVzSpDw646v2+LuA/rsLSCb/qbySU
xJd6ZFfdXX1kzJfd/DBcH6VrDAoFY7pgRYyCzR/BJcHWG16/3dpx43U0iVml+bDoWpADcZ8Vrf1D
7+OFDv8QMfvGHkxLou6XH+zP/r4tPGKpdiy84utD2Du99QGuAgn4GiUlakIodHZ4qDJkT6/23BnW
neVBjBjhi4s/QM68kLDDD8Dtooj8WGEvIAkn7dtrS1bf44ICin8ULS18WcguzNQkEeQe38+WmUIX
ncubRHVGSKH97SX+Ak5BVIYOdVsQzXs0HTC9SRkpPZqL0pqY64i7LeDa0NMeeoOcTF0fcx4f1+4K
JCHzc6BsYCZqNcHkdYnCPCYiEucuwWvfhxQ1KBM9s4JDSP5YRmPGsQnZOwtIDlL15EQ7pFW4MoPr
K9HWTyq8F6ZZS5pVaez2UpXcUnDcc0kPbazq1GCjAeE39zfssPGJPKyDQBgG2Y3msxrfhsvGIMsj
c17rYlertYVVaNDIZ21TaXPvFk8PA5am+Zodsnc3VZDwsx+4nOUhxStVz0vbJOMrr0+ykLRZLW5t
1qVn5oPvfNcokQVAlHh1O8lja9lRHxdnoNK/yssg9oJ4ll7UxA20Y/72vshpMvycd5HrkJUdvyNO
Wa1i1p9fbMUk1NA8HNI26UuSbuq5nUw93SqzHs6Y4k8cUpjTR6IWFj7GzTQmd7OBy/hoJWtrqhKj
7OB5SsJza8Tu1P7RYr1Ml3ZUJYbFqW57pDT0zB/8CCcrw6fe211d2WT8UXwOezlGfiNtoyjJX4co
i9jzJGJH2fROgMGJDntjsSsjU4uwGF+0wNJXHeb9olUrdGKo+7gj1zZS25Na06BXGNRTsexDlyRp
nPduHYa8g9Ar03yOde69eBkT9KmnZLALRzixZZLz4FVS3s/uHjFIjYIF+takLVEGcA8NM5Ft7yow
57jqrxiafuWzX5wB2XesGKdI3iaoet9VdLtu9ZbunwBT81f8gGgeVoJNXVIFvUckL+vsYR6pnhVu
NqIxZlS+TDGdvdysE2c+ZhQVScX+KuMeCxtWzz3/3rBE1fsQ/+YqoYFQ5bNKFj99UUhysiANBo88
+feqT0Hr1p66MbYTmCIsywv08RAxrRURiogv3IFkKCYx+2yOAIbmNTE8NTKGDdMeEOK4L4Tm5lH/
5dBQAgQskCChSoyUU8GUwADODHpZXoXCW8swA92VI1/3gh3xhNxNRtQbzQaDrTOcD/wTnu3HOdN4
32RK2hzZWgf2Vz3yU6Uk2HvnRn9YIr3TAHde81WCiaPjdcxVwsYZmH+QcRUfLMSCRQvTwP5cKKXZ
Mf5VjT9PFDWLEeWQS1Fo3OTQ+PUrvGKaN4ufUnEOBIzJ3zGTX39z+7WDDr4XFJUcV7cQ3RNU362u
bOidK/lkAKHvv15R3Uy26wDUcQif5rvTrjNgDzt77nnZoShtW/118adZFiI4+e/JqzE8D4LMtTWA
wSRSCykewP2kcLO6aqk2q5zTbjXgAMkDz/hQK3i9rmsuBsJ3nvfV0SzFUtL97TjcwdskIw9iAH0n
gloPhZkC55T/omPLFoeI4EK0e1tDBlgk7gnYrDgEqg3SAjnhH6c2K5W0NrqZ8U3d65GgBpowr+Tu
735iHq7rovRrOurWeRVY/YvyMIPDUrUfoONrS5jZjzAL2BP3iXTS0VFqI7nyhlhmRYWLLmVYsL+t
Jz2zSDxGVpgdlDvFUMHSpFYddiL3DJk/zvrb1LrIByxnTcjEPrLdMqmnT6rsBwjW7QoBnQOWN/bG
Fpe1XhL98pEHfA3YPplceVw3luyYs0qO55lcaEw7qcrkJXLlhWw0mJ8RdiVZoyvFp4Mv+MgwSPnb
J/3nB1TZAx3Xme+X9j/N1v9Nyw9pY8pYcrfWdswg4LgVZveMNK5i1RamqGCUDlfv/kIcbn/zNrbe
DyfGKHlH9ZNbYY+E2c238Kx82yWOWCdABGwlAKc/HxsNUB+Rl7TcPhnRq20GCSNwroPDq6iQybCS
RXVEqu3kKKkWW0maly+Ls2IN2wOnnJAuFZmGMe33NoeG7RZUq2wfPUrU/lSY+BfpL/CdmF2a0Cpg
lnW5N+tOI/f9VbbWhP1yv7is5ABLaHNykNmKdsbfcO34yJPcwLr/GhUqhK5AQLDyaqdzZSh+OXd8
W2Z7AcM/pNO9HeM+h+RPm66tfL8+M1dUi2Nt9XcR5N6cdTIQEe9JYdtvAkKVzttHBRzf8tWoebft
mWt/xQtPNqSWT3VT0yYzXiaq2t6iTZlkaHru6Upv5CuiJAGQ7bU+Te3updlgzvU6VxeIBy77XtkR
BGs4b9/KP1ATY2y38mZ21G/qeeun2JE+KUafqIRsfl7BlvI5Epe6EMzgEkKJlREzlkLBbfPbKdk3
Hntx3ouPgW9fkgeamCiKEMXp/tNeGZNys2wXHJgCGp2BckAVqPy7AKGgtDR5v5c+my/TLkeivqE1
rzXzAfaz2q73ttq3WH+tKOO3q+Z/IxNmwZey7EKgR6+yKAGK6PrNvRFL5+DUt1hRr6+A2v4HHgr1
wpyBxuu7CW/Kwswjhv2Me0oso8XF4v1JEpxU3F75u5ats06dnQyrMBRBejqlPKosHdYW7+0Lr9Fi
I46eyjHP5KnW5S6V87mRXH8oBsZX63YPvsIZFIJ1cDyPlBuzfU5BjjtfQGMdPlInRjdAyLJBULC6
svNwCTLJzgRmW0hp1o/KbZDjcu2MVL/mPqo2Fkb5MGI3KCN7R/94yOu9I6pj/jXPkUlIUQqEdRiD
OuJR0HNzRZKndU+X1jU1Y23AbYXyuHlEV9bOyIOn1jrwPxy8hCwImMgIdwBM+3cZHQPAvaRF5YbD
Kb1i4Kpep+X67hCGjczwAk93gTGvvdqiVzNEi5iavFcajvqbCkh17wjcilY6xzPQluYdtkhp+hDp
yIaIRlQ5sQzSQf/2AQF3Mbkzi+2sOsOzwsXO8pUOuGlPC1ToHoNt/f5gIS6nejOE/B21tDEybbF/
u9rF5nzR/RfDshHd4fChnQ9Hy/NTIQlko/CMYUZnscwVqAZnvkhC0D1ktZ29f/Vf6lovDENcBEGi
5uJLUCW/GwqVQQpTnLsCZZR09DdW7iicEDvmzkJrl1w0a7xiCTsOKhcygqcIoaODYkkLcXvohdlT
5CPAh2qXl/Xm5tfewAAO1Hp0sxaNWf/u76NkAQTTPEmwN1zgB1pS2J3nuqNnwqYypdffpFtjqSoH
Q36Q5/y47XvOqGa4sgZ3zOH1qMC9dH/MEq1q2hj9gKozhVNkR6lDhfPRR9KNvUSHjGU1TjiOkAgj
yxKgstutripIYnn1QVy7hEf8LAfXqk1RT7kbVG/ZcMZyszUYx5kUG6eqDFzn+9EuXfISc8CpOORM
GiOkcVIQjUr9dX18/8wxYMhOZDdI/DQv1lk+IcpM5Xs7R91PglWl1fPj25Kvu7m+YA9O7H1S/rdi
zfIPt+m3zCQcxACIRG5jbDac3f+hw9vnX5tKjHoYr4jVNYe76K+lngcSPA3Pil5oofE3dblfT4nK
n3OADX/YCwTw0suemUQF0co3zl7++mgUXy84P3GA1tM3nkFWGrSiAcl63wQGNkhK6P7OPKoLlWGE
AJ+DV2PpGRYS3Z9tz934aGkqApxWn5bwdS1RI4MeS2uPvNlNWhpJe7ZHj1ThkPiscJ4UqkONzrFz
aT+XQz7AMwFRpYWp0iO9C113jUVcfpyP/SleM9cglw0llv94YzENyzBoMHE/juqqQH2FYsA06QUX
aFVGI18hlEFaKrNxGaECftDNUukRWwlOaVCvbLnXO+RS0kv/YUQTRlbUbTBV7JCga/3F3ASFAmHV
jcwr3+0e2xeC+qdeh8wIofnfrJnFJIZDy+gK0iZ2DeToG4+B5Fhicr335pp6Wk6yYvDc8fY07zYr
0Y4OQ2Mgp229M3OfwuuLQ5v9HRMz+Sdp3Z+cqkA7q18Vd60pthjioOfcj0t2epobgmsy1Tm6zU/2
fhSdwmlWZ2me8M9BYhVpYnWv9EijSz3MNBsuqKgXh+shFvMdREdWJSA+w1HkgHbmtOewnx++5SdO
7WKaKoADZ+jGGdCsI9yhNEC2grWORi7m5B6foRjJRd7Br21a/NeYepcewZfd37Ol2FFhfqPV3aDw
A62tOyQR7usrXJ7NttVPgE+IKXEBLcynPf9cSFMORWyTMlcE4QKMZxCX1115Y+hzis9ub2Kbtrlr
vW6z6wzvG4gdczLZMirU/EW3Q+GbVkM4bMrgyM5yRIfK9k65et7A7Wr/3HnrM8iWktLwt+XdDcIj
KvK1mDFI3nRdNHMKeid59iDISKVDeGzQJeZEH7qjxbmaEQoh3eMxw4L6PFn4w6aCrh4WwawHAiCr
X07sIC0Y4hRMOO+FseRbkWi7AVXNUT8zBSeiv/6lBtmDJcIBRaNGrOzhpWxg6+7Vzp3aHD0C8Hmt
ssUVgiElt5QPgsWOxpRFY01QZuTGvoAk8nupfxx2eGNe5idOYmGD64h9Opc4bTcL4GdwYszXS4dt
KBTX/y99iK3q80KL9afFkjhYXUFrKNhl+WbyXMzygydndUnENf2VE8lL7pNuz0uzOsTZZTZLGgWz
bhAhbK5CHNcIekr/MgvrGH3aYh5djtUDRSkh9nr4Jb35pIrmoTDr5N38MfNBRFwQGAc34zgOQbaf
cE/JRswHVqcyrBU3dMQXYhkVrhsB3/wHXSu+DDQ+BqVJtnMF4qpUGIKmPzzs1IacWZsJF2jQM7pX
C6FiEOFLVEpp84kKcxkXtoeBHDACniYDwvr4lquVg3754q3xaLalGn6sW1l3zbfZ7jE+TQ8enftg
zP8tJ85147Psaeq5TYLZMybZQYymDUtfS7PSVxggx3aHo8ifELPEP146aeiS1BeYHUDZrtc1fgxE
tgxEOlT16AcxTM+e212L0V+QyHUMfh2IPYtzF8ByK1byXdYJ5qA0TnqS6TeJaJSZHpX10p8SWQ/l
PrKHupxCbQxcYgJ53hzAc9FZLaxH9N95CX99D8Mj34JJTeZEHfSgTwM1l+cmitSRt5MAeousw6i+
MJcMTPcvu2u7iZbdeX/Vf1maGtGpHLTT7k/Ihcc0+i83S3xLBl9PddZbSwVwqhf1CC0q3ZsWusj/
v+5YodiLIvyfHtEyq07peEXuHeCIkBKYrd7bTbptX4kEIvziVUjXLUL6srywsdj2eMDFcuVrHON0
E7JiDJHo8oXbLYkyztlEgaO8K3kSTiEhOIAUCmki2a+KSdXHhTLtCFlmX9XhFa4CdN2gEEjh1XcL
CzxkIs0umyoru8pI5/rX1We9rGqK8UQ9laz+vNttx1jgj8XdVXwoOtF5rxeBl2umzkeXMwBQqiQb
iefSLeoQmub2hwxAt68KLHKyK70Dp5IeRsT3Nj2Rytoer4lcgEeQNfr2yUX6cKmg90S0Mn5Fnanl
SFhi1Sp6YvJfhRnHCbK4T6ln0+mhzwh+Q5JY8qUnLRysMNqTVMFY1IuM8FxKD3v2ggUS7ngWkhBf
iyLQPA7oL9WcIOA+p4JUwV+cDqXFClUi1NPUfsWAUat3KiXgxL/QG9i/XYMRibYXZ99DHz2pBcpi
2E6gowSvIwmwr5y7JK6IB5uxhkfHjqedu6yPpgDi8Ohhqm3p7fMLiTSUlBuATvgFhGKbgB5Q5nMG
iya20ZNkGM/+KGZcfcQne7CfkXl5opIkX/zSfX/IHHlSxqe635dBqS/Qjd+BYe1VaF8c39diqXwP
8rj3aq9jnemafZAYNA8cKptUG1BKTFwg7NygBhmQDi/PLyGdCtm7pA2HVWhI4QHPLmoChptRZ+mX
JRhbTSVCRh53qwWjkd0Re6LfNq5UJ52HBtwxOUFDUkxXTuLbRj4S9L1dXuIceV6ZwVxDJhZdihkD
WutNpxw/sCK2w7/AuCIlNsdT1qq68CARUwZW0c8MpcEDZPK8F/3Dvr9CO3KqKtDPLYYWH/xpTEdi
FHQDKmpIxpZeVAy9QkfObhpHaGb+7GRu+7prDMkYEzaGzW4fh9hyu9UMoHTU6d3e+Rs7/VYjSrtb
fXVONzoU/i5xib6TgUDw4Q0ljIdDVKXF9iSSxZH97JrERa9Sgc4F5FA7KXJmOUjx8+DrIUVok7sX
C0BXnN0YlXiozN+yNfN25AaQLlXQXr/f26A9usxr24Otn+I2aTyWJtFrpOafHmex3Ef7ezIIZUwe
/qXBt3l7XyGacwN0twobMygczxaTRjOb/kWu9oKmFi8fCCfLK0tlMjEatO+VS3LiRLcq1NjCdmP2
NBBlhahew6AmZy6xglOoFQ+QpJai1SIORUlA1FXnFuujvK5BM4SyWVZfJKOaDOdF+njNpILAii6g
7EydcYJ/wYkQyx+0YmTI+MeAwKQA8iawvFWSa0BIa1I4t7/HMCNBWjFt1y6v8rYOSGS57fvhcOiD
+TDzjHFNSApIDE5pjGijG2gSgESenL5EOgiMOsQFRn2vBkv3/3D1xYA3b/P0c7HSaHfa3aEFnuB0
zmtUmpj+b3AmzL1VXazVBOjCBoVZKW0/JgrYzEpSIBjMyprMLTVu75EwVav8Gf7U7/AK5QduwTw1
K2jquVSw2FgwonMm65ia+BjIC5R+O8UQItqnVaNM3FIc6VK8BEf+tzo1g3uxPRywERNFBc8l7139
KGB3YmNkaF+vNpc9t1uCa51gbIUdtMkltQD4JPtumXSdTUurBjlTo1FgRRjaOfzOyUvA/IYISzH/
zjbNcJjzWrc6quyJAUi6KjPfXzXF9oI6kBFLuw6uAaWipxMIYxqEcI9v0vLIVuSOoLh19ugxpmuq
NX3iW1WQxtcU6EgHsEnsx5x3mJhc3iDirdAlee0fjVdutsY7gZGyLvzbgRf5O2NpNb/t+uOSxAGg
ea3PBYQxcJuAr7rSMt5JwiPW+sc21DzXUOpl7wGf7u7n+OQ3MgL5qj0Bpt2oTQMx1jaJlR2z456r
ay/bfStQMCx9u9GU1yX8U/s+uedHRVYXrRTPKPlfmtVHfJtc3f0mOe6ROLpWKTeLlJ9UI1vvi3Uh
A46RyqZz+v40ho0fWogH9DBcl7T4cQBZ+rr6Imy3+CbaAgcIcHUt38UHW+lp1PQewFqRtBB1cCuq
PNTMtHT4Ad2wOpKw1vQ1jWHeKTi2l1tWizvvPvm1YcFItDRhSYCpjUJQNrA0coYfeiAdCpG56T9Z
dlJbkYmjAKT5NBwH64wp7V3N5r0/GYcElBw7BcfDfM6wq+mwj6fAg/zI/Yg8ii+gnlagaDMva9hK
QxTnGo/A24hQrF37/8cmFcE/HwDCXn59zEBViEPdyxkMIIk+H+m3mo5GChPt/eubzOoe3dYT5riw
qJ7So8Slld4QL6gCceD1nz/58zFyyF7Ng+pLYyAmq+rmLMNJ06FxLxZBDQ42RP+a2Xs2yhH8Xl8N
htjmrN2suIN7aGQ1UApVrSCfilNVYa1ObxX2V+9v5LtSk4GrKICyJjuWo7Ut19BCyPz+spDTAIRm
joOLlEKoKTsf/l66omigfIrEH5pQeS87boktXhwbaLPQiSWVP2AaqNrV+vd/5kkLbCNTEqFRF+/g
O1FEdPa5Sfydzq78gWQPa48CXX0ITq/2sNPxvlODMlzBGMifHbMKNzLl/YTBXW5g9HtppM5El8gr
71olO5E7lWaGhpRMECZUFw7aSlb+vyDM54W+O+LVRqQzURqNOyq0h+wKBUG52J7dGDCWImpRWTZ/
86vOvjP0mDVVBuqJtdSsPnD4vB3XECB0CvSVvac2CaJ0QJSwKg/DOJCvtWSZOIEreTD2UoWBuTTZ
tjd+w2knpbOVptcDmbsbppcGY3GowfDmDWsRYLr1/8bsHYCeNOCdve7X7YDALL2dsxbwzOyDW8om
m0mRERbhRX/d0DinWpmUVMze2kO/FZ1CpJmFYGqzDeALH0u5iX0pY2EEdLv2IKG4WAJqUYcErRwF
irHAn9NjTPBHoDWvlMlx/5FFX5JYaZUgUKVGp2i1oxdQoF1bcYIwkHYy/AuJXHyhVrfY+QjYtvWP
wymc30Ex6bxZLJMDK26ONf31qbSkGoqOCjKzpC3X75/NWXU2cI2IAX2ZuR7euOlhGW3kGBmFT5kY
pfj7Axo6lYEl01ULW/Zr14sfPtU4u7Xoyx3Mdos9g2Z4tz3WwiYoJC5uj16sN1vwDHkgav+O2hpe
aAAsFtSdIy6txXsM/2ew5qbK/m5hjK/6kEDKG1e0ropPQuZ7cKhZPs56F/xtZ1pi4+qkKJsbtaBb
azBPtd3gRNKWkEj0z468PnvjJ+asBaY6Ex2LcfImkRmhvrzKtgOxOAAjdITLF4ZoZYjjBUyrPkBx
HEXflXJt77CgBPOcHuE5aoCHtLUwZRktdIK54sMZnBMQox08cMiYYMJFziPklH7sEk1gxvMNkh8l
yq0gw66BsTFvM2goutNccWcpuKUo8I2e8xk20I18pU0W4UIZaEvzsiyQklsO7IbiI5RS4G7QHH1x
tiA1P2IU3AYrDs03Xsz7TaZ7puHeavCND2V3MleKVSlmsO3h73PJtbmZ62b62fPKgF/EP4GaGZDj
j/YqXlwL1ISm2V8Dv/2eEiWmDlt2piw3oyOtIr8hCRjkUT6+hJDWaifriosdVHJGF/NalU9/n2Qq
wyLfnig9BtNHwwvurJ4t8SE8WN1/TtcW0hNF2uwtWMFW0amcye1I1p3mWtvD4KuaxbjHYE1QmDrG
Cie+PZu5HOsTYdmKW8ofYXQoZGNk969FstefAjm4nQsesNULJEIcYgxUuhLM0Nhd6LujcLdYTEc0
JKtGYf9QwSW+a5qApVxMwuLWyau7sxQjeJgIi4idWom742uOWIi89eyp9+kaWp+VA6y/iSqc/h6I
DcsVbokDepqCsBPIOuRS0KqEUHRKgD87yxaYWQSvvxTtwVE1KbNYz4tf3NVQlf7pBm14cOi1IXyT
FKML41IDuNT7/c8+qhYRrK2a3lAjbmzZWOA5PhLwjkmEysykWYuxAa8uBgXlOuRPPtnb7PB3ghT+
s4i6Pht1BbFU4h9Pbjqz0VkZoshu3Ia13X4kVuA6Jg8OPEEt0RDnXRIwmAz47XNZHM5DJ9vNjQ7O
b6n1DKr+AlMVhBYPOEtoW9QxuHIzEb6bxcJoU30BYTjfU3SlymYckPLJaGcVNdHyEK3tFLJxLr3O
h3vw2Kgkxo5jMChEFFvfzovf1/lpqdavBqmjK+HA89rYsDKaAKYX1bNRwOb07e13qbZ9iaMNLPe1
uOjj8ZttXtyVFe3Mqdhxu95+Gn7gAxXrmk65nxXXEGICLhvxs45LpVQuhph0PcW6ZBNavCLxqrju
rfxVNpsxmTJ5FEytT76KMb0HBQLacnAHobkxzo6+OBXgqVPuUguhASNLNiYzz06fqEfp0s+zczDP
6jKyxrIYUBD6eVtjkrnfan1W07RmNUxPWE6jI3xPktYVwhIuFNtLFuHAHaEC+A1jHmG8uTPDkKI8
/WbDMHv4PLxqqegonTpflRkud1QnMlrIADAb8MtBVxraPi/weJqi3e5mWEcwRujAb2qesMRvWnPN
s4Cotk8PUY1CHc54zHx1mokSAI7xLc/HJ/7bLGXXwj1SJ7PDxEtqneehgblfU0gVlZ0Tc5mT1SO+
Fl/dlVrgFP7JYTIfiNGusgFg/X+T9Evx28hEFhgDX4F6/rxjxyJr8CGkRwjzCRu7w49925p5wqtE
6X08+El5Ao5sksZbEp+DFOLtObjzWkE21C6r99Hu4RZ5eU7zO0u8/CFyYvSYmUc02JO77HeF7L1Q
5U9+bKzWV63f0ZbAxHqJkw5GSoxOHixkqaT0y88RqogbgtW1ieomP4a5LsG9N7hLUk4SRHptSfbP
YB6XRrQgtb8XQO1aIduNi9cn0djHhbYmPRszb57RPPX1UgZvheOBVnOjMA3My1XRxCV0N09Db17y
fs7JtO7WQB5VG+V0wyLlGWLMcouMB/09IBsZxUgsiKknPYfv/YQ0Fs7TwfcAO8g1TA7li6dPFxuk
7f0JWECL2CHQnScGUHwXYCqVOiQUHeKppq3f1v4uvdrjTx/eqY5T74QU4jUeyixIdtM843exbB9p
OGgqxAxfpBXZeJxDjY0+qaW3gUmi1no8jbrBTYLsYptVFomqvURpmGpEHFkKMEjsYgqsJ9aUknQ7
8hjYFvCc1Zd+Qtoz9llRy2glYKQ+iNUXwz44upvKBPp4QkQuMLuXb1H/kwvhasPSUd86SR/1wkWY
42VW1FSp9D9MAWWY+3OVTgzP85eeN4k/UUcHR8YckrYSzcXHDrSGeJXlGJzKPi/nE7ux07XLXEww
xe1Xpuhb3aH5kk7arNKFXk5QCXHa9SRI0usvDGfcbblqVbIdEI2jz4CwWkyF8Bv6Ms9a6Wc0lk93
PLBPzeqqokSclvASQJYxyA29lzelo2jsx1kqC4YyUM/NIIRkxVuYOfwQyPsC6l4m3Cd/8DBOLp81
gum7XBl/lXG+yCpBTrxr1pgZYZXKWRNKlBoM5Ed6P6P2YKMPRY/KQNAOcntZWhTEINJsIoDyyfa9
EJGmiYx8z52ykkqn72NrzG84Zdy7SBiSxUynnTMNrvO0MiBZASkXfmSASo7JzR1C1SAHZv8iXmCs
lhm7M2xJ2DerLU11c3rNkhlqSQZ3YHYmV6JX+ACXzwkG5IH8OYfX5XxClDJ1MKQjCVeHkmUvqj4R
y7He9aPr8o7Viiok0UbQae6IfwZ9rtH3ALQzpUKb2i5X11MDpboJ3YDUKq6vkabKbG4YDaoV/u0W
B0/DL0T4p6rwlli/53FiohJhapgXVZjDzBroKCpqkDtwEtNd3nl7Linn0kM70n05fqbmp8UGKtvX
BzH8YYkVgT2Ky53tZNyhsf7RBnpfO/SA3gO7Vwz0cqWc3HqfSBYjYMI1aooql0JfzS0xJ25PBSuN
YCAJBPMdQDTvEl0REvKhbzyuAzwf0JQLg+yIALxkZac64MvySfLDGwv5R4FekDI4l/TuKw+lEBC/
ncBkZOsPFROmVZhNFqhHclHx7voBBApwnEKAFqIcDzFiB7LsNsbtq15PJIbd5gn3+l7tB2RZFjle
/KZvUrUd+ZFFO8A3GREcr/5E3/LCWPuMvK0IDbe679o4S4u13x5EsuMefaIlC0d6CEy4qswse5ge
c3hB+zH6Lg/8vWCu8T8JYpXkuK/qNGZiSl4Lfk69SVM+maI5wvywl622rl5io5z/BtJZgGQUS1TA
f949CAzYE9jBCIxlu1GDB7DU8Ws4YuMGOZmq1KwfEmDZaIQEKQhPUK8w/duVqN4Z+JAih/rtbtKz
F/8FNag+xVFl5J7cXXRgHLLHYYaFPCjS85O09Khv92KjILGrcCm2u/kLZA2MBJDdYIjOsInOZpbY
EZHKgWEaXyqdljG29LfX3/zaDaUhJR1nMe3Mon49w5nLi7AWbTz1G8lCQv+Ll35G8Ny8AwCrcmnr
Tidg07PsBeawHTglZjO2h5B3lfG24RrVRYTX0NXr+qpgQfB/iqCFkXawtp2K5MjmcA/tfFX2N/2n
tVl2xc0kDlasoxNskPUi0UTVQLYXuK5qoynlz1WrA+QkSVDlOIW7IzvEf6MeCMy4VMo+w/Fw5fcQ
0DCduDI5pn+ZxX0Nfg5u4RDBqf3yIn4bQKE5v3F31wZ86/U55WY0+WVKz4f9AhO2B7sfPngHIPZA
HZvjhF7MccsJVdFSbLUXhoIQNJla6vSfB64rJuxtGdDvzL8xUd0CYZ3bIKNsz3r5xrFaL6X90QlF
9b4TBcLsPi5/uEvN+INC0KbeFE7Oep0epP0fSKGtN++zF0k9ucCV2oKeeVoX+HJP+ROz33EQpToP
TEREzkCLGGfZFy/pPzY5nZQeft+cBUigHDCq7Cywnz6qSimkwrt3w9g1NAq26i2le9/ud2p2z8x0
wrMbZ8xISaiCk5Wshc4qvJKBDEyzmnnoMnYrtNtUWVFs1Hutd8T2JDF2IKt5zvFet/PKFg624QBf
BgXuCSngrSG5n+ByxXlGRlesUvt4bVOLMmX6e66v2dAi5z74wM4/1jLfa4fyrW27Igc/A105Q8Kk
CNIZemdHZgnpluKEjxQENvhs84mfsjToCjlcaLAuJX+MSnz7RIAbSXTM0KHRvWeMMYCfbGdCa1TV
3z9vSJq5lAXd1duM51j+h0/DlS7w/Of+dVkSvR/rd17KUwAgnM91UM5JduNb7pj+zUTA1xuErOvC
BzgcaAS/61drhj7/vNwdfzVPh9GDNAcMTLtBwGbb9EwR0JGOmjMCXHDlQGeefU7XpsOgv1VZmCa7
6P0Oa8Xj8CTwMesszbP/cYdJ8nJOXEnFFc7fTcqhjPLrBISr8hOw3PvBQHnkEAgUH4vt7vRAWGtR
ynzOnQwRF49+HLS7D3HHAAjH/A5ir7XLRdgMbL52ZPzSh7YliiY2V80cNgZKI1Qh0uXccyPFE2ji
OrAK6BUBKt82lXGXED23O5ZPe1dP+5jWmqqibQf0WwmTBBTfyXuiDhAqtTLoiWM4NuRmXYtnQpnZ
Z0SRD6kSDFeC5O7xYQtGI5bFy68ZoaKVfd+0IVDC2DWFF5CFPxkOobjMOIOBlwAGzdTUl4TrrDyE
ZywL+7i3jZVpNpWAc93R3z47EJ6P5w1bec0Y4Dq3Z1HgsHFoNg8sDc3C9ttvyQuR/ewSUPxX2kwz
qeF/QAQKLXM9WbsDN6E69pkIwYY7LJBVcVJCQLc/KvBdKERsBlzy+9Qtl4nQrJVIhBa2MNczXIU9
Z0w1QmRGRo1zENjkJeVld2xtIdNMc2z1G72GDW/jMv8Y0xQuf1BBASddAF/3NtXmKebs4AK6t1PM
6WLKPKMUdWk5+kccJVnes7Uo4CR+py/vz2LH4U//Zhu+X2s/8AXlXKl8a26xg0Lzvipa9UeGmnvP
chWJPjFtm5FH0cnGkbdb9gK06+w1XlmSgUky30+asgxF0zbWDqgtNn2YJ3xGSpFlWbAiNA5t36BL
xPGKWEN9UByWULhrCO8u/CMiFXCvS2wTfV33YaBU+SI/3qCjXBw0eNxKJVnZ+MbshBiFA+31V7pO
3zqVbpnz542XbAVet6/sYWsrQQtpOpg1sSnVBMKAIsvfZdMen5+6Up2W/sGFK7NPw+03yOT1Evcd
w9gHV64O6nj8yuNoTJk8eJD2jcc+R0Dq6IfJgG/b0PhuqDL5tOjn7GzubOVRIDraGcmJcFfyTgqn
T+/A3/QSbnjcwHuhmVwpcbpz3xb+nr+DjvpQg1SRygZCOxaycGx0eUu+HJ9iNFpqbmTZFVB3127G
manYShKhVLEktjXvojKsks2qqPTfegDDOnrRq12TkrGk9/AGv09xs17P/j+9PMav7fwVd3gJGiny
1K3/WDdg87q9mayHap21dDowbyx/ekwHerPV5Cc1dua5uiZcKEu9oyHRPggpjYIzw5oBFjQD59Pm
Sy2n7QByCr+185HKMCdi+O+kq/TcovSFAx+hStEWTgUpkdOWHESytXMEIqZRoTI3DfYyZbEjeZC8
zXNqbSxgWWtG3OV2TrT2D2X2/t60VqC1ftDu/x9VcZSbKJCJG4lrZDdr9TLpR5PFKP2CAKo2UU4l
A2ewCn27uVVxYNX9MTs29wO6v1+8ZZvW/9gFKdmlzLgVTyqJ6unEHlqrvAx2AKO2NX8nHLvwFMxb
OUIFLu/Y/+7JRNDU5ENpV2PEmGtLK+uP8Ts+e2YC8+G4OW29/0nSULbbEdkf8aiC+rVeAd/Qx4+Q
aZ/wezdCQtqV37RynA9DBIJv85x4tXDrgMz837d5DxyJQCTunsRxF5ob+uz+lrOs3wieU9Z7EKBd
11KD5S+2LRXe8Aohs1JApry+JmkWrJ7gABLm55Ks778ao2xgNeJPhL6lseQAhmKnFCO6XjA1yegd
J9trEHhoK3vVsFeZ9jTMpXTuNObWa61b3EK7dV7oy+veN3ovHrZPNGfn2Qnbyc5+Xl9muE4b0PQa
PR+06PVBmfekKvN8qACClcdgE2tKLm3F7hHW0NHK51RzJgf4LuMbrGUkXJ/naaNRiMGyf3r95tn9
ksPNlDkc1RifbkY4GpT2b2SPZvurRun6khILHLGAyjH8VZubS2XrQr7Yx5cu+6ZKRP6PKhxSe3HR
htSjCJWk6mFvJsgLMhSFrzZTI0NjNL/rTkAfUcR2EX0/WVZJJTzRk6JLELmxoFsaLGHpUe6r83x9
DKO6poBIX2G6Bqhnd8Bsi7UNhCreX8TJsazhCiACeiqzK12N0oJKprH2O3MVRRKQkYyVdnHvl2zz
CJRtvyXyijTDJuuwZXq/0Z9T6XYWHGcgtFKiZmHovBVSCL3c85LJ3Zptx+h1J/FeziGyB3fJSA15
Q5wNjzyoymNgrdfL5ArTwX0lBp2OfT0GJqD29SBDjr84w5zvq3onD0CMCjBHybL3JO+/lCODgb8g
y8D480z/AMKRGg3rflUdTopR/EZndxUEcmYmRdJa1OpOIvchtBtFcISk3hR5EMQjkZiFbdTw+Ulo
FrSd+GQWEl0IPhUIdOlD5CQObW2Xuwjd+B7bfcZzP8pXO8MFDzAFlyeFQlcBDWKeVzb5VhqoYkPq
fylEraortPcM5sIrqGBBPpj1J2rAi1swKKV77ciDqmF2Ybx6iSlu6soJb6wIMAPoKz4KLfYHFIV3
WZXNUq+Rs4smkjRIkH+xNMjdis1elsTTvTKIE3ephawhkVsOs2lfRp9udsTxNI7Xc+hOv6igZqO/
wZup3VstEKRR7r3ttz/9K82gAgFZfVWoco1pQjnOSt+xkcrTFnrAdXNKaGAqGQDKUe4vDtd2lx4d
pTHrqZUUa1705khemeKvh3KMV/D/uwEmll7aKRdFEvOcIRsstIzDH1/7iVUdrlPXBBi1/U0/oHh/
FSf4X+aOpJ6DfnSkpeFBEE8zH8OK+5X1+r2T/1L+SlGvlH8U7qp+6+VJuCT/7P+E+dM/qnhV1huT
2rj23eHn9GXaenlRCduBIDkxi5dy0s4gZN8nb3sf2S98itown3DInyinFwOxqAaEghFjotIZNZny
pITVrKzBj+sGx3zc2hc0HwLExZO1Psw0XEzbBtBt2JyQB0y9pn+6Mh6XSdBn+TvNbiucH5TQnyya
ao/Su0cp5CoocslWlmTmiJzX9XSj0c/RVx5FI8xi3uv/DahTsQ3KxHitJy+y8LB82TZQQngQyz7m
D+SiPZTPrwmB/OshcHjvvHcfTMB5ZxEcKNGpAyB/hhxoILgk99JrFF5miPoXqSS6ohstqsrBQBz5
axNzJpfjQ+1+XZ8YFs7LLwJ5O2Hgkhjr3RJR+HYp8mJCNrS7BBICjAe0/TvSf1ODKca5KNcmRdGB
0LUL47ApZrf0XpQl3TvD1c5srx8kMJYR8kiKO3J2h/9zZc/I+JWYEMUtfMfOV+ZgzasB9RysAS+E
OZ5pSIM7/MYRC7S3jzF5Z6jwvE5XY7deYOQ1sJL2FiYgyU1/HhTNeksIGM5kyEz0sNgnZT+jAiJx
CXscdhHMw33O6pbxFnXkZzCDNvkGd7Y+uUN9BeXg/DleFg3CrAWIYr+2scsMXaZ8ZrLMegsj1K71
ovEkQF7w/GCHMphMO34+2vOMwpes7ZUYP4DUaejTkudEQKGD3CXeAAn1LIecM/hdmaqZShzKF8di
HRbvH9Fe5Mf9zekFgtmrR07vbPCUaQjmaKZjqE9SUW8v1bvPzI3axvSv1vq4m6pQWlyMp7+ikhKt
lSMBPKARsbZUDYtSzyGdIFf2KLrxiwHhhru1ZsFpQW5w5k9Nk2dryC3uushdmzgF6ROp35dp/+LF
hagFs74lQAyEilvr+FjjbrvZn5pqlkUum3AEHAqk0Xhmyzc32pQn+qTc2KyE4ePsOk/9cxzPJRlG
mkxtL8yHLGXnat5mpAotGldrU5CjKLfmxZLFGJwzxQquU+HoABdMmpaZDr8z4mx/vdy4tILWpKcN
/mZsfM1EnDRXQFXbh0QHgIn6EsiT9OZYORav6hFJD/d+Cu+Vq6MB+RQCFBjSo6ihU+3umjo//CeL
BTVMYX9XnP5SxWLwm62+ckBfHWb8QkTsTJtGELGxO3JlWeH5oj0cE4nOdm5n057nLdnblmKj+Ww+
F3qtSzZtrFhirLdC/KD+aVyZxHYK0CxL0E3jjxsaiLG6dc/IVDUawtYmNDhEnjcPQfhV5PHJQW0T
KgA/H2I2mo99hz4V7Q83NeLwma3FYZ5FwV4DKlg/PAfHvTRpd/sp8oJ90udaOugXMgraTBnfhJyb
JG4brwLVVwg4oNpFeRbC8RVuv92wEcnrIBTLXeI4YTMeyV24N/8DDsBFIrhGPRjI1bNJ9dHDzbAn
2Ex7DucxoVioTDEnJadfOzQEnUyfwEjrYVytcyvcdCnWj4vZFV/YVsFqurqNRjTNC3KMG3tDDOQ1
NxY3Zh2VfPfYVIw/dRq3XPUxLPMcTHE98d9GOUvxgXyKarvDWNwFqEdhFyraD9XTEbbBoKfmkmxl
StBIM96kXCsXUI2Wela6zCoazr6Yn+Z/DfXMTyWFLYLoWAGbKr6pTHBiR4S3Z8hXDox38Zb4ezNo
D8Chk4CHxEAOKJCerW7iovawCk/I61rF2drXh0yFmkDuSztVHLjsdlUcU8a8azr1gBL+QTY/7fiD
6DpnZiUcYIJ3gKy5vURdEfbrR0TCeEj7BA2K7behwb5cjYKZXZk9UAVXfNnm0Q7xEChkWTf7J1HE
UoLvS4DiQc7JeQIIMMDhJqYEYpzS3BfFAh5RbIQxfr6f13szf5EkmUPKN+8g9JDSpCcMv6i6FinY
gPZaoSU+w9TogX3PPEqwtUUU+C7G0Pz4OQse6bvmnAwpL2gvPMkfBW9+dlYb1WxPfBv8/kEh77LR
fMWPhBmBCvJsjqqPiXD8B4evcqFZrS4Rs/VV3sE2vrFzr4rbEnUmeyERbyXqTWXdj4xzBczUnOuZ
OPUkk/WL/p0sfKYLldDhY0Kx18Ga49YLX8E6AOwahTNAhMpTXOI/2na37d1FWrtFOwiF2vzEcid6
9Zw5m1zrJmKFSnEgbvDodJ+pQwyf2hZq5MXeqFTfIsTrbnAkDkbAYBc6kBR3KXddw26+Ni3moT/r
/xzIaAeE5NBFAJEz7s0GhFrEBQAZvGZrI2E5DgBr6sUjB9aTFC9tIXx3l2rziZXMfxSFJEKihZQk
ZfQMEu1Aw0hVcwN4dITixKbeVWyDTqb7GEjr297SbdP/Wkdy6+GvpaFryRr0VF5VYaL2V63fGhdx
y8kylTj6IjQvzUclT+K70y4La4vhNKv7N9vGCsodzwxXSO8ohXoKMY/Xj0B1j25KlNMSglxVr9Bn
xuYjPX/ePEJvK9S/NRdu4clKOZ1d1LOP8sTieyePbcIXA6rFm2AhV8m3Eh04FlYLHpWQGARIP/yo
eWlIQm1xY1o0ReC7CPAi+lOg6+bTi9N79JXxKValf2BaBZ7NfBxHJWRB9JZuwcgkjRY2ejT8zW2G
AjaPu3Tm5F1qMI8UC9WFEWaW3aMXJnlcXGi6c6QApkLcuRyICl0VyMCLmdkQ3WThZaGoR+kklODK
JKzxc9GAmCcvLQL+kLvR8v85Ohu/2eHN8EvG1K6/WrKo8gov3P4DlV67jLzaAJk7Vho9n+XueT3a
wVYWvf0en/FC9HC6jjqkEqZC+77uRZ4ruZafnirU7idZRa6H/JvRHfITgnn7fwk/uVStY/dEh7Fb
szoMUbU/cUxiQyDl/Cz4dmLjd6D2M/zj0eJgsTCZMjnworCcGJxfNgm8fILetL9SeEhpkMFtovXJ
PFkwCts7/ChtZyWObvLPKevFZWWjW6aK835JFIae3NY21nfFVwLNIVk46nUl5jr1xg3P8kyQcgJa
Nc0SDi+iOyBms7XzVcrcV08rs4B2aDN5y+TKqQDJD6/mowpm5JIwwz5aVORKVQsPGYxEeF1scEej
baHO+O2UfHIHUOAG3NwTdmLravwn4mjO/O9Q2gzaE8X4S4pp6/G/5Ge5daOyRHZn6f3KOxOr68XC
hm03WzuHnKPeLYG6ZXLF7Jga1xUMndfftUwWhyC6JoJwCM/jBdmmCPB5llhLa5MgVWMcZLp+ocg2
/x2on2C4OConRKff3y85Uw4sYS/2u140VoYOsQZ5a96uDpC7VCVKfhtOOTJ+5hzgelWATsM+Sl11
ZRsY+tsvhcv/XMImZsn/DGXE9DRCI25ESZKMP0lo8YePZt6Wk3UvI3CugiDAgcptTD+qDqdx+Ixa
s9iT6MKaHcU5PSe02Mo7YwqzLVpeQ61FOTfKnGP5KQvvv4zB0Kp1ucO+c9WRB7+N55VWEzmQpYs+
6imlBF5v5tVDb9qb/9NpeIBn3fGfpOVLe6Bml9UV6QR0o/xxSYPC7RAASkHPSa0kW5CwWPr2FqWC
nYvJw7L0BC3mXOCVqezoH1w92WoVOKi8HjyQgp/4CybAr71g9ln+bsJLk7BibTpUQVasPRTiYXIp
EW/DgxnFDsHmppveQVXhaYd8Ncsxve+YQFNdaQRdmeUWMF1Xp0rgjqSyzxZ9O5zj/FCeEGbvxmUt
ilYn0AqRXiqf2q75VkLRdkuV7zHq5iOa4JjtH7Krk2+J3HQVn5v481/yCJtFA5YF4/ZvhVJReTTP
4TdpINKn9DrPoZeZLOVRyxgLuhrCnzsVl6LGma+YivmjyxbBjwJpyTznssZcqpAdS9g02CTpB09E
vgZ4KyYpCK0avWzLZZEjHuiNq2xY81Rs5LpTyw0Xf5f8ct5HdwHoC1G3DH24zmvHXz/hbMjaE1GH
hRyT8v/LNJqiP5UYbRc03DgGg9fbNID90+xsAZUFx3xw2YNk6/ZMBiw+elZJGJXUb9rBOfhkrKbw
CRReshVJCVQlWJvicsFEsaSA6uVKhI9RKK8oRDrxloDrW9lTjEOWTT6vKObeMZNfwUfkfM5+Bkvi
/pAPgRX66JKROWqjIfSw9pHQNyjzwktBlQ9yeQ+7WpmKkiHN68Nv5GoRqM/teCjQdQAyxsT8LZ8U
8VRjhGgUF/uiNMiLKab0Va1v6Z9tHuc1XFfOrD/X3mgG+IL9/tNBFt8tqtTpDEieCmZAmcObBrH9
XQj3u9Rc7rB3E97qzr1uP+qqvPKlagFAOM0Rw8N0wCKxSkaWLw6TQUu6Ogvg9f7RiN8eKbl7+Br6
Z9Xv3I/X2CHsAwUd0c9R5O0fIrRuV9TwEn0WQuki0WeKe7+15+epP5JopVjSj9uUIMCJrxYM/Rl/
HOqL4Z+oP4IOk7ITxYoTroJkDLltmRFqsJIhDXfw7ALJ8uzYDfD/s/xOXBojgPd20GL+U/BxgJSM
G7oz7S3Ip9n8qDFbhNZrMKSLYeAW3AS6vL2FVLuPod9UPCnTtYl8zztVj8KUZ541EEZbDL3stJVI
+0gRlHM8UMhB1hYiFTRf/P93bz2/xcouRmmlFdbGVF1JRiRpt+AevnnbWICfT4tXQuVJIaHP8rlx
q9z4cu3TFrssA2HJDUm+gm0gU+Gb6XgNWK9WPtG3fUkV9fshvpUiZ/mHV4EEHH+zKQMEREuTIpwO
IfKGh1WzChqM/14DKS9N+lkfKLO2uPOPMz/iYyqDaBIZ0EahBqV0bDTOlTcVi8lryoNcxsVcA3Ac
Jazt/WP8GP1vfMVmnjYaKuOE8MfOrwCTJrSoo5eg4z8wRyQOTaQ5Dn9yENBMn6F/5G4CJRhapXoY
B5v1uOOOskexREquN8X4SsRYbwaH+Nh6sbOA9mktkvakAxX/fRyxshxRNz+MJpD2DO1xKNHujjvW
b+F2OAP9QSS042ZDMBXwazhtRRcUUcpuMUmOZBBT+qdSna1MkDMw1sh3tNCXrPwZccts1Tk9zYyM
Ydm1WKgP5fYbXKnfVkZz77a1pUyRZ8dAT/ov7wpIJuNdPh2P5/PkCYXvkdS+9v9e5HGfGFNroV15
aRIrVIZ/SmWz/SEjAfRzqVWjGoHUlpALWWBBWvC+7C2OTPIbc6sT59w8g5ev+SvEH70luptnzggx
mXkJShMVpEjWmk9bme1Cuw+8KSjSknz90XLcNjoWOCRVNKiFi2eGLu2OAJ/Cjm92vpHmntzBmcMJ
v+TNYx1GfoUfVlTYzi1kQEmIIuNPlET6wDWY0Bwej93cr3kFiFRtC9lYKA0WVX4UB83xXaBK12dL
Z/koQme2kaWFd1lt58n25yJ+VTTy58vorKiw8HQTjhOxviJf8YwmJfR9sNjd+7YIuYp5CNovZETt
+NIMd/gBVDbCvHniA//KgMT1cq2snEczbP2b6mpkPPKW6CVSu14FXceRAnc6k2iOAqmDu/akPM3G
LNISVlaxlqqkB1tSXRhD59f4W4BIEijU2APqRbEuZE9xm0qBhq5mL11T0gxQ0HuerR7ca1yNseEj
gZd0HG2fr5cX1JMRoT+03B0CCUzTEnaB2nfewacuicAchyrgWsEkS5TOir3qdI98uPDeYVR19Apo
JbWsUs+2REU4J102papVlJ/DePf93g0f0bD/HXMJMQn3GTz0JQ6dexlqY2183hvJYzmXvyOkAzpm
pnyPxAse0Yhvt7+MS246sfkDrOsdu989M2E+yXi43GZZ+x+dq4h085EreD3/zNMgMA6okfL/pCTo
l5/3D9Kob4oHNgzDVqdHO0wmuJ1Es7plH0WFUO7vrTcFCamOO3W7O+S6X8DTuW23DF8EMNYFOlnK
cqhoCtOYDGWsFiRxvL3OfZQ/bKILVJRpBgqixhoKcbB/i7SC44cf2w/mReNfl+Srht8jAnoHJo7F
UQXW4USfomuHBFkWaAm3jv3DQyqankc6G8aK6NTqNmuZpLIicJNreXhWnWFmdNLA8nD+qhid2qbX
rKuDoXK3SyovK9xBXWM5RL5U5lrsF6z2yzUeQDUFTaTIBJ4YyFSWcDKx/AupbRNZpN4UxxCbxQ8K
XwwbEVJ7YhLE6D7pdyMJpuJ9dEKK1+m2lSPPCuLRzm3YYC0rAaa76x+5O1FY0yZGp1shZKHPLWPt
BhI48/Dnji5o00MibnRGflNTS1v2+dMVZj4WuO0S6wI/LSdS9fPVJMAyYqamtlJ0G7+S2BTtfpLN
7DSrFUtN9yMWZISwfGPR08GAhvaoMdEQj8Yvjple0Yvj20m9ZVXIelZY+cJfXOHdc/BXaBkOAcz9
jUdgCSSaLKfk/xKmbKlya7UuvnWxKEbPyfRct89zOZeF2905EvTPFSluKNiAHab0A+xY1/Z3MFa7
GqT/VvLS/XBtBswZ4po75n0HvoIByYG4pRCAeG6YDxHSU+KQYtKYwYdjhjPu86m+pJxot0cTgZkz
5yE/RNs1Kel+OBru7wcnBGfUa14s98GB8jXnD1zHIszGJAUsg929Ut51xFhcdze8a23TPPqxtIYO
oXQM1L+8E3XihGe7KV2H02iFSs2T9mj4Bms82K5YqakQq8zZoUdqWubAQjzrlHgSqMcgLo7FOned
lsQpLOcLg9o7b0RMeTpp9udijrXfPzGl3L6KacwLoPosPd1U/ODdyBHg5XQAmaDzo1W0XbtN0IWZ
7hcq2eOO4w3pkx18vBLaMVwGgN97/HrlDHUber3P3TD4t0Y3ZJ2oZSC8DflaQhTTH8YbSBuIY6gq
5vNCgOvQs8sP4WW8xyRLuaPQIFZxYBszOYuJnkqhGyRWkdt6zKSyel00vVsX5JDJCVS3iAuJrdY4
g9dhBAd4kn+56/x5vAv614iZO+0rFVvnhStYXuGQjHY0vojoLHLc2dcGEYC5hGKCrTV5T57ndY2G
hXQtKQdBiuNsbh6vFZ+HKiWZ6ga+pZ0XQ28WDprhvwTFbDnYCmTK0Bxz8pdwzdkI4L89brVuXcIO
bZqFBubuzAZY27CtKl0Bi6H7TZkwBGlHvcbIF84mi/aYW66gyS76HO9S5kkn0a1Omf2fF67+69ae
6s5HGVcyhGg6tOhKH8+eig2ajj37A6nFaqimYITlgxk+C6fFTQt491hZ2Q8XkdsCRyWdH1bCD22a
wDAxwTglqM0I0uRhgDsOh9LlD0Ly9nsAwNa0WJqKAGaCokdJaBkXucjn45jYXyjSdv/YGYHTpSvA
RGJGnz8qetMRucrud3joFQC+EdbVLc3g/XjUywm+IuYGUlAxodkweusTGU4MwCNbGt8E6n7VYDMs
PxuQYeI7y+okfRUBJ9i/X14TzKK1iY2Rw/hN/4ouByRXsIpVguGL5M38XprC/F9gVgK3ie91Yl51
f9gI3JCB3POdfZIxH+mN7jJeBdBzIUsdh76YgGsQAPmvHHq1n7nnhUo7mFP4jalaXSIG5P7/K15M
5RjdICpTfFU9duPY0lpdtsLvuaQ7jhN0V97DuSjkzEhK59GjrSb69B3+jasjdss1GhnfPD/Tu9pY
nUJpa/e/C6IocaKzDri/5YWZo1oOiMMRXi0qxsOf410DdYonOV6QBtPGUunwHsq9BEINQeRpgurF
OEL5NBd/pfdojrq547oEPVjVauJPvmzSB3aeODSjpHio+J1ZGUUSfTFnUSF+9M75u9RhrBHdhn7c
Rbqm+kVxuW7rfGY2QyaAMf4l45iLwVoyKdjKQ3ZP48Ok1MxqDuAwZDG7aBPmpnQgfge/17tiKraP
u297ABFBGkEZtX6hvZFkA2lnh2Mz4fH6NBHWcumWvbsu9mwR2qodc/ZJGqE6FN8g9Uw6uaG17e22
xGXnqliooMZ8mZRF1Cenv0F6ts9tn5uwEn0U7AdIAS98yWEnpWplPgaQvLeNE1IljS9KbhRITuia
T3vLJ5XJhIYDhzPsfTfq8sfd0mDkGo5HSMETM2y2kl08cvLaTwk3v08PmKOsmA4FoGE/q0vGaUVt
xcygMuAHuoY8Cepxf7KqIrFUb1IKvrxGEN7bX/SWfu48DDV7DTak/N4bWvwGO4deUdaBZi4K9Msh
f6oVVLkoCe8YuvKWnHOrNw6PDRzzkxnT6pTczxsAwnm2Xmw/EEv+kggLGfUE5fBkbHweEznf2a6o
NhAnEpxh1ZOoxedFjmZcShzy2QeTjhr1/FS++j7J4Zl1R8XM1Df7+7kGfgdRbclsytiJGn2dyXM1
5a7asmKc7j90zfr6OA38YL0W+WLh5QZCcM40j+PJko6PigUGmDTkokuDdQRrhfKvS3iWK2FL3bCH
cvBxwAmgyNyuhy2e3P8wvbXlfgLLIS+EgsutofWIPwD+qjOKyrUR5wF4DlQUKzJUI9Jlk+5Wd8f6
3DH21j/J9u+H6cm3Uv1IwgUzgqSX7/sTDgrdTF1eX5dGUp3rW+BaiyB05h0WQuXNHjXDvd7x599B
BcDJr6RBSG8hHYFMlUqKmorM47yZfHwS2yLh+dUFL6OEA2e+sXFpyIO/DeJCQ8AZRaCSml1WKR+P
IeZQJuwlqO2RapdAsRR30aR5MbqokSJNHNlT5rKwqKnYRjIftY/Hhpt+7qn8i8XIdg2aoYnNLqAV
dVOg38kAyQ0RLq0E9H4LkT+E19ZkCNqoMRcsADOcxVYJnWJBZhyI46Sonpmi69tQN+vEcRle5E0P
3pEcqvE13eX9YKjjWeBgneKuPScFYYTP8NS0L+DxxhzFHzrSvdQv7PurR/sMK5EUU0rX+lYx6oLn
vfWjjLFgKeIY0GgzCjgAWNEfAKnWmdIEPREpz7NM1QNV7bSuCk5MZEC7Hsv16Mrkm1BuQAikaRWa
3IqLKPPAcUo3hiBQShGWA0sJlLKE/beK92umZ+3qNHR4gaYlhYv/cp7uFUq3VA4edxG2+RTpRVii
2bPVy/nalGaeLtyoILTsSBSfCV5CQU+3096neTav+aOP4G+p0yXECEriOqsyb76KNWqe2KXUrm+D
1gQNdgUHKFo+/KsFbg4FqDtYI3PLnJuWzPP0m/TWmErWfbH1sQmtLgBYzzYQ/uFrtCqzYmk2/aHl
MtPIgbLmeep/aTOg773ewt/K8ZGH7bhr3eOZaeW0nRGl5KYzm+ri/olAYzQeyj3feuHrHKPB7St8
4SWPo3cIiQR2WMsIdQdEHzfDgz7tPtntbADkVoGy+6LhkCM38OFLjv7yRmpUPIISlCISGYCPloN9
sUTZyCBXfKF7avdreQyDFxCAYJDng2Gb/of5sCaMkjO22WwRDWLHmTYyVTT6gxfF93RS3UVMPtft
e4KaVy697GSjXrF4shMIIop0ffTCtxbg/ePGf1jGqhkWp0HFkFqYLznPzCPUQLrYNiMVHSD0+KA3
r85H1inH1aIbPm4EzW51Zeym2FtiwrHfjZlhAKxKTA1jcLLEIxtkO0KOuoB3xPpETNf+g3TI09vY
vW6f6xaLwWKYUoqx1fOCwEWUZntMobOkdWTILP34HITvXqhhKquRavlgPZLyW5ObCsp3OmrAOF3p
GgbsUV/uPqu0Qdgo4peHwXosJ8v1ehAbllfKXWT+NM8Zi0Gb4oKV0V31GExaFb7DvNCEibK2VYBv
sFwuwZbFiw9cRQLmYpmMvJAJqy+7xgMEW2QIv1H3W1TWUSN0hQAFPbqhvuSnbcMUBByz/moCpJmL
VgGJlX4gBTmfQ3/+lAmEdBemCHpcQWzCJL35CYVmeGEMUlA0iftIeCLodoHdHHaOUwHF2Fqi1y0i
6n7MhENuAKhbro046nsV/Uiqc4KE8/i+alwAam6dxwjdH1dF8BTk0FQjF7s4k+wgPrKbyuCBCWRt
Ij9zy8LdOJORBkrpO1llibZ3pYLed9rrR2b22YYPgpOrSR62RG+SiHB6oOzmkCo6eVZifJIz7cZI
kIq8gZzgdpi8MoJlYZ04HvldaW04ZZorCkymIt4OiCmAbV706ciP0+rFwuTRjv/4vGFCGf9WUR85
utlrh/BbUKhVKXHi+wEIy2GsbEhdNOokUDamRh1FNuWg5kd+9obizV+/4seNTmVKSPzROKxPQskK
1/Fdo2huAvNI2b0V96bm4LtwSOL8M0sHJAMQ+04tT5LeqNLZ06cPP5jcuSZeup+4yiJIRXD8JLHc
zRvXjC9drj5ziRsd7eSz8nCp9Z+z9HZoNnKncgAwNmkYLwcjBtTNLOHD8Zvy0rns6bXzkT32pTgQ
favml6Q6lYOlrLj9B9TKFxSzuGniGt5StA/P3eR2YjK0iyQ3Z643fKaT6HEh4yJ8vgWxuajYZ28U
wP1E3+Z1bfrKxe5+hq0WlcLGj2K4qIFKcS0eQIbWgUAGQAx2LUDHx6rexqxzvtDMgbl0TkMnZ6BP
5jMvPFDmB+FJkojPFrHzt0Cl1WYDC6zhYOEMLRAe1oLx5LhQMyRPNuHkKstCerBM1eGsBlwwxLMi
GaFoDhhRW33nRd3Jib0PqLjpg3392uoJC8EfKCWd+AbjXwd4s5HEr758RkZ3WKuq8comOVd5YloK
yBXmoQqwzDp2d8Xo4lgWUmqc4U6zhHGtxp/dPAOha+30DmzGznc53bcswBVhAFvM7eEF6ICsf16h
KZNRxQTBX/fCoXpHt0Y8K33jznwftrhmefq4U/HB0keqYYmrRzsZFhmjK9aJgnZUINAXItslbwwy
upyLPDkuL0ax10e1dAsCrooa5TF4GOVSaiYdvwemw61mmVb4o1w9z66n/UgIedcj9bg7tpbFfFhZ
VuREDO9pE5dM3tjSa4Wm5i8zAUD9gzkbK+fpNzjblwUJ6v8RzFX+TIlcchk5U2s8LtamoQg/006Z
s2P1UXWinho1LQSGlddYI9i0mwZqzJxJ2sGwJ7k0y5Gi15qLL/QPpoen/h27ygn6RRGy4RTRUdTe
rscMtbkNc/dKxAsqp7BblqaraAmSYYhcG7+liIwwjr88ujk8o7gjW2cJ3KQjWFOBohHQioCfz/hB
8coZoqRWZSh+PMAwhO41rUEW9iCJTFDYRp4DT5Q4SJzF+CfQ8dsLeQ9a3gQhavjxhXyjcwu7SHUT
Zhrd6y7GV2pPdDCS2aPOxfkwikIgyT4Xm5XdjUgpvDNX8mXXllpWK57quzg4JFOTwohxF3wip8Ux
q1eINwjEhMBdrJo/FjysqN9TWkzi4HU82ySFJmlSQYIxC5LdtD/pYrSyK57GCxRBHsgF3TbFpfWa
OvD7nIPYqwpR83Z3E5GbsUcCjCekh4iNpc+h9u5IuxVAR+yykMaEF2OH7XHjuXiUUSPdD2JsEbyV
JJzBqDGLBW1No2NIetkPX+v3TImzBxMCvPcs1TIQZqmUGgV00UlVQRVU+eTLnLW76eiH7TizQlur
1o54Gn5LlTD3XHMUc0gInxZDBRgZ6zbSpLqZLEbtt0FYmVKNYaYtOFFyMHrMsNfF0lV3D59QlofY
HabCMsd28UfyU89PFSVeFTQ1uifswCxwDuBxYzPBnGENLHLOVn67WoQL+XFchyIFvarB8hQnDhXM
79q5u7nVdTxUoLISbFZJBIdyuhU/gY+9Twsz/17esl+/P/RYqH/cgRcLYeVmK7a9JF/2CFSsdBCN
UNnp+HPCpKcJFzw5gMtXk+Gl91Va+WUMfXZHJ/GiDawdorMmC3ymGxn7FTtNXckucQ0iqU/QyJu6
Cp2Gp9ttJp3FBm/YVOvBVAkxyTl6oCb3GeYNL0OQLRj0cLEhzex/xawFLQII2N7bVNk356QQWPYR
thzszi/XWXeiQ+GCDimX5F+MsgU3w3x1kFS91e+opvuOZ0ka1q0QP3EciufHpBH7O1bMDIS+l7RC
vdaBub7FMJlWzgjROfOnGuHAFCdXlYybyabOBEBb46C5wD7/dIS0JjucN07AYKxGwihf53tpDnBP
5V0itoRgVJhHaHkDwWV86ZS9X+Tcx4Ck8H6BCpokO7sk7tRGTxfJ3RPw960plfTaoGffx+r2ytZA
s7JzQjqSjbGNUiv3QqzGX8eDQbxuaM92r0MZdXHalVPOIUbcb+eHrIcq77fGVraK0hlkrWA9REnQ
DClGnqOYz6sRfsYQBdZLJxwW8rgD8rqGidJoden5WawLtQXkjm83S4hda9xdVnTl8BZkJCXO4RGo
qIR7NA4CLCMpJioi/b5Q1cPdHFRr3MeT255484HphN+rYa2x13JzBwsTV1WT3ThwR4gsMSowPobc
y+cikGDse85knCGtBZ2Z3bEeoCkvvMC5DWqrT8U24h8/x5FuvN0oEAEB6ANnTcRwqivUiHj7c1VZ
rR4p5y8+uDNL/n1EjvsE2hsbE8H0EHQG7wbBXp74ch2EoPPggGsQ6bBJPyTuL7yPatX5MCcMz6Hl
WCHbbKikuAVjoWmvu9ZAK3FHgFUL/ECgW815zoQOFv1nAspTviE8bOV2YCoVKzZVR0b95RA6xzAS
BYpUXEq18Gxl7mYAFebAkY0s/sYMM6f2Q6TVURJMuvn6+9f/1K69Fa3aKsWYCdCIyl7zp1UwGSuX
ebAqf8PbbVdKnVLa9yxLXoNbUvaqi8Vy6RR7zMw5UWeV0PptEiVvTB+dnDEW3ftX5mAhCfFBsLCs
+zMRuno++A9GTnbOy5T7GpEwjav02pPGB3QFgn7MT4RAIiaOfUZkdYesEcootaoswshFIJl4s/XE
J73P/QIFYRG/ldP0LeqxgQ0zyWj4Jm8hhg1Qw8+vVsLKAuvLkzkYncOfjcV5EjczBkhC0GmYpmHz
X5Z0mGksc0FOFbOsldh2MAmPG2ly4CDR3dqbceFs2LIFdu0B96XkeBV9U/SAxyVGB4xhlYN6NDy7
2FjHar9A7ZeFu6wTUAwaVjcVRX5chVfKgF9gIQAZg4c1N2FfrtcWOHK7u6x0rdyE/W+j+w5w15CT
+N1Chkf6WE9ZE9v/tiFt/qHFMSqijYfmjIgXX++oWdI/VcMsGNdNpbKbbswU5qxwgCUPf43y9ACq
ETf2sfrMcvRBtYi17ASggoPruos/qSkQksPL52WI5DBQVNDNQcA6x5gOXE8rH5eRGslWdxshtWQG
Ww5TmxDXRaATayaptEnaZMlTZdYiVZHmzEKJpLLmCaCYZT0JtziiZ2LD/s9c3vw9biI0Zssvygzz
kf1jxypUf+reKM3LiaFZU+HG2E+M7v+WMosyZvQ1wxQqirK2fzUzVkDa2Tkr87c+XO3avegw+4wv
Q7sgli6Oz7VBq+IkoS3UjLz0PWDRYQ/So4WQPzGVFTiVCL6bPSHGqYLCmP9+k7CH4bWO3GnQ7F+a
D84NZkpHNzZ5M3BIIYOLH7PuX00C7RWXn8qOvHsRxtnwmupmuUA5hmdSyCR9SvjYDGlna9g51rt8
DHP8p8gTf/S10A5n/ZYmGUiP5hiBytuQcE+w5JdgTnhyXTMTVc7xBoolUNnU0oChDSUA/54b+b2p
2ra968ZWSDGeCrW30BTihXIAdVt2/6aNlbLgm0Eba1zGqd4GjDDk1WTMpVQZPc0TLqZcYHL7A6EZ
SEJ+MAXqMnRQO400wIPzulY5h/YKHIDW+pQcG5fUb1/VVkqNtW3682QaAiMeZF4M9gSVBk6OrYj1
1j70vT3/LFYZuUtoxswZloHO2v3mImPbQ6tJijv58Gnw6+hu0b1Si14Pl2/YgIMrmiA45iTnw5Om
sScMUiqVbGLLwM9taH6Ac1dojz9nXGMGCdJ4JJrJxmexEnhJrlq5qX3dNeQAYnjciPG5S8NdH9ud
EYoWzONN3l9nplYG1eUEn51BxP5EXC0W9/zOnyp/oAdO1xLhbMfYBDEH8ohXAR5FUHV95S9POYcx
OFntSQZLx3tGVZIXyNLSJSgRO+UtmCIOHCl+5jovf+fwBceWkEgJefCXHb2yFgtpu7C8VxG2x9XA
5y87n4u1AnKUDpXzZTGm2gsasEMo9JAqPL6RCk/Hkin3G1vYZz4AqL4oJD8CCMvmaRovZNaB+J2/
d0pVOoLjxrQ1KBM5zz8rNEEh6CTNNn+b1/TaplT9mWUBIqCouH5kc8FKCB6ZTR6csB7JV2uBJBpV
3SjaFZe0L9noxIQ1WT4/whahmBWmNkH94dQvrGEtyQKW+9J84P//v1DlkkuaOrAdhJBitf4cJPRS
2pjt7DBtWpUsDKwGOJu2toPOWywnpzqrheKN7AXQaB05O9TVdEgyrI8TY/maCXQJ2rlYevCkh07F
i0IZGjR6y+jXNv5g+bAPbnPVVZurzAxsUpxMm2OvHK26tfjCthS4m4RdkZRZkxuFxD8D7wiILmB9
00eib/JKelMms6nc6GTWow1GDrXizZ0AO4x5pyUpD6kaGefo052OKeaBrb57IjM440crt2JkBSY4
+aY1BoOTJzxpLfeMdQRp/E44uwNs+KIC3HHigqBcrEVAFDWL4azksloBZbtEvtzknuBEIcoe85m1
FR2o9mJY4V86mry6YTpZgviJPvMMm/2OSnr6MUghTra+IsrWTFfC4fqUep6OBR6aKIR9o6mGJDOT
Xl/vuSeF57aHmHwPuPNFF7VLxeAY8iNpibgCIskpwDmhxKAT6zxPxIGLtay9+mm6zLtMZLatz00l
FPRWf4qUHD89oRxoo4AVFr8aZAavtLuHCRvAp957f2z4MtD3n+MglzU2Bo6Ewvzsy/Odd0sy191u
klMgTyzw7BMQMeWPgCmhYaCh/aHfVusg3AtZFqexZFPvb8RN0yqOtVGhGZtPRDpfTv+MIMBIdZP4
wLV5SsItFkMZxPdNmUz3Gz0xWyvzK4+FMQL8NoRhgvm3MAVH6cUQElNN6ltB0YXp9qjXx7Ha856X
bgw2T3lX8J2ktWd0uHybd37y3IxfDvAHWJAmS5hZZ0uUbEJ0Gb4tk7GpRx+K/u6TrJbfH5T/0AtQ
AV7CF+R/nvI/Ir/psDjYOtKqzZVxk/NBrvTNTNJpT/7RaSGwyNBhNiYy7lzOOqXa2ITez1NOqTap
Yq07W7e9GXqxIpfps399duBfBlX+soNu5KDx/ASR+thO8ESu/2ZcWib9uoMtBcZdI40H2n/f8M31
4AUSt8FCCLs5d7lVsovZ5THicFy93VKOxDsf79Iwn/USyeWOfnHWY7NxdW2lKvV8NcKuK34pXuzI
wu53k32nFoQy5pdZ+gy4WJHRI9hGoSZ/82TwrwUwXy074PbixWXfL76Xeby5ok2rkOP9cZJKvkXS
5HrkGclvB9X/sTSrewTiBwwVCklZHFZpL62av8XvnCUzU0R9cGM+kZo4lw8C5AlqvgtGGFu6ch2y
LapyWhWBrCjERm1lbcHzoChwuZg/JG/KeVFoqNDhuS+99b7DW6isC0agCO0Uenuj2kpuCC/04yro
q3ynxxw/nQbVZsFxU9lKUIF7OP++77VNeSzr8BQgfkgpIc3zlKLTRJWBbY9l7c7e3+KI0zEkNAB9
foowUdiqsvdAmb4iBdPxa9fuVg8wnC0zAlXinr1Oz2/YFNrUQvFzTVsq6wi6Xp70+jPcPudPryOE
Qd+wdsgAPTp3XuoB8BLbjOHbvel2jgkVbpqxLoKwvHnFZi7dY2HzlVbYO4zPFYBXTeM8mHVm/0l8
i81GNyVScXxIeQt2StAIa/oSjmkCYkZAWoBkErm2KP0FuTQJGSjVR7/MVqg5R7P2GVXMTUhktEqJ
Mtp+S6cvkxl0S4Ek04g/nJyrnKMqznHQcIQo0CqV+bZqo55GwtRJUwjnQ9j4njQC6FSdmossgb5R
2b7ocQ0wY1/8vFi93h+HUs9IGy3KQ5R//c0jXBnrly2HCFOMEIBKx/5ca0yhQ0Dz5c+Nr162kj2w
OuZKYjVLaI7fHgfNqMzinpAtOcqIPvAXJa0AF2BU1PRpZSIo/wPgoSKmXwLoLDvFVPflTlx7XCSp
TOSjSL5ii7Ho0L3mUu/C6o4ySjiHc2GdmPlwMfx1SazpZ3xWLVrR4l/YLT9b0MKvZlm1uakc+q6k
jm1gclwhFkBWDcLMPvnH94Bl/fbaEMDaA23iHClJYgEjyDEHCO7k+FWX3J3Cbxs6881vvUL19XbO
9DN4nYmh/zMMAhcDsg1ZHgF0gsvIGFesb6FWvu6tF5ClEIWUTs5c9wxP8OP3V6wqOEQAZ052nycD
yXh+ZUolJ+CLfikP7Zi5vE2Ig8hVRlVgTSxTnJgYV1XaQdoWGDWMkof1I4SbzRMeq/fZQKGn5LjI
HCEhzaZ40gHjoQExPLZIB9OSjc3aMCMQ2Pc00C8ij80bU70mNw+igY0N7E5wWRlpuDtYu7TqKO/p
BUT8os9bCJSVtniHhryRQrQ2yTT4H+E/nNOs8zJAXQ79jnXwNJEUgrNNYQlhk8KGEL0PcKpOjgSV
wM9s8RLw2gwH1h83lhH/qqZH1GLVtHFA2smqJjqBJc2/y4i9ByVSm3C6dcHLrPU4K/6qLz9pNEG8
lB9s/4WMWtb+Br942eMrF0c6IOP2QEAB0AXHg2UnLOdfObRtmlql8jOj4BS6EWeIy2UORgU2ZphS
tsu+CfOFf0amQWnJhKoQVJ5lUikSsh0QxbA8YhJlvCUhCDw/EXIE8z45kBEHNhlNA5C88oGWbbVz
tITbR/D86Kq1u1Eq3268TzPgOq8HoOGbKJhrLk8VW5qkzDkbSjLdzlxBXZc+5CXFJoX2DIa3kRA/
ujBkU69swyuyWhXm+pyryfkXzW6LoTG9jPfbbH4971B0Ix8ka1T82xE1FGL60somhPRwQ5UdOY6Y
T3JkaFWRH8zmDLyHqVj1L21yJD50UVIrtg7eMsf1I4pPeltNY+3mYbt1zFAjXNebG4r4Tnh7d7pq
L+1XOWzg6uSHorg0x9ocNYtCH+QcXgPJdVe9FE6uXtRkl87yRhFtI76BnbkrQkAEfoxydr15LXUK
0RupaolLsqw9bWSMzbJZGOZskHI5HtpmN5eTQtWt8DMB64k2O2I+U5JNs0wcZHA3eZN0gFe6ASXR
IbKK2nQa5ThbaxFcdGjBbO/MgxHFpJ6Dp9jmjSQrqou8jvFKNKbiXVLQS7TuStF5SuKLKgKFR8tG
HS76EjNxSIKFHetfQRRIP2f30trPG0Peq3C5043b1KZsi274AP/WtaofAl1dSxlfujdRFSwV4+DA
8qsU0AuJChRKl6orxLChPAafLXHNC8hKTy6If392/VFt2hAOPkUnKwUCPmy9Wuo/+tWWL6GaOh4r
kWiOTExEccOKPR6VsbyVzp4oocn/D5Gquno4azFNsnRZpFgE6XdiGuw4bQWocOUs3WNogVE9gAIQ
5UTBAAf94fNbTdsi1D8SgzMpL+ZB4DlHTZWeiWlPaCPM1yTJwyclRPXq8+yNo3vKB9wxYC8Foqfm
EyAYG6lYLKxc00V2L2BG1fQPLLIOPjyiTYVClnb7YKROTIrhaPsweWOFTvnR+zJCnHqlros+JGwf
1ihtvnvn60+9504ECklc/zjJewH5rNjBDbd7KjBH/gKUfk9sq+b0Ui6s8J7EbUl6IvBm7mPVr+Np
yO7W3OBS+Ge8hbx6wjHt7d9pdWr1L95tdwUKGdkc1d1UBXcO9hgsnXG3OeJQeMZZ6Uz7JbXi3b3U
cStQE3Ce5Q54488g6PU7sSTjcqnYSWD18gH4V1pp4hI0Vfbc3cU4Q9/lE1Q0HVfROgWgRWFhgJ2v
NSS9hoREZ94cxsHSc5aGg0Jv+xusR5RTLWmciBruNbURhOl8P/VfvbTwA+KQryLd3eBQRVJBfI+x
WC3Mi7XXa7ED/9+h7aj9K94pqUuhWfXMLmb48q9Q2Q1qb9S5B6x8x23IzCh+ebuCwL3dUKArs45b
S7jN75a7JQ4jPhPXMW6PY4XlyLkB/6vrG980aTcs+TluEkOKlfFXTtPo98MPJLmJsqA+QvxQtlXr
zl38TTsCUpZIVl/J85miyaDFT5WhmsCiuRNClqIAr/wBBlg1ISMDp7MieuqRFJRiZCfeb1ndZSH1
JCftD4wM+Fm72rSSx5rknODeD0eZYgFClHjTQjsgoNcICiX1LfplHN1G0TGZbuU4uwcUNNqcnvR8
AiQJoMsNmxARGQltTS5eNnaRDta4Ttty8YFdfoXIJQNXf5g1axW6zkxZjPCono0c1a55nTcNVPG8
QKRwJujD0FNus1kBYAicGxa+wWO3AUwG+2ExRozr9BtV9C7I+Dwej7TBfFsC1KXgPCUlqv7CVOWA
zRjEgUqRW0KadX5g5PMiy+vpo5vW1k0E7C3i7k765cn8BbFsr3AYdMYK/0t+Ma130oE0DtddoevF
RFrMoAISIRcivJ3JaDhErJKbppDzHWOH3rflO8O3gybABU1Z0cgyWPH64Muj9Od61QT2v8HdCzzN
yXpEadVS1FEB3jW0Fl0QqTO1RC/EaveCaGo7nprrC3+M8T6PnDJXHZUjcO7i46vKzEWpaTXnVk2L
9HmmDu5ax5ZokfA/VOe4z/FO/CVB3MGp8G16gMjELwrnCTO1jbtaek2RTffWmC/EisT9yRZfHW3Q
KtbHiPZb1D+JyINQlHbQh+E8ZF3CuGOCzdf7N0nfwSnzVSkATJY9+TBlpFmToWfUqyhCHygklvVQ
NrBF40ZOiQD3+m8e7gTlOiIPDS0VqUAvbU1DyeNTiDIYO86p38ZFnEMPOai9cXXEDP5vTtlaiAGe
M/mou28lSOVbZLgy6iNdFLEMeoifskxvo4eaWS7KPFTS0zm1H6fgzkxmRTi05iVst34MiX56lQs9
2GdrG3pZx7fwVM4lzA1Bk64CFqpNE7B7dMV4Iv8UbyHzKOEoGQigfQyZ0noxNVHXnIR8hsT4uiX1
fk3UH1IMeHtkIsghUBdqJnNcIVv+sUZlKNtLlE4YASjoCe/ycLvwSHAVwz1txRfsf8B1L3rDrkGX
+idz8+gAyVEBL8vgX+Ii2WYeOpM4BT9D6hnOuybD3gI0G6cujBsWoul2QtUq+UW1umCcvfvXvsPX
g5wyY5EH2IbhaMSemQkHUo1WVzxa6dldWeNQG4pjPK4Djlcx9O/ijVu6ibQLL52Ok4r25IWfkPfE
5FbqDxlCAo+V9T/Ak3h49YTf/COLdxVEXzbyfYf1jYKOLpSxg9vCcH5GtcTKPfB83gzdAzZFJSaS
qpQB68cPVnsVOeN7wg7At/bNeNPzOeXCxcnzoRyoy355f3791/ZTyDdEwYQRnFX88IvxD70CqKiB
KX0AvMghNsPaLR5KEslmq8cWmpUd8mNkHDJ/v5theLFhTv5eciO/m7sPFBHlVjF33FiVpET1sxmY
BuseiIzjjssb27zCHzVV0GvTfdSruTRzK10KrSpLYIAR8Jc50mWu8y9IxAbAq3C7+GpYp7lR5387
oNL4n7Zs1I9v9CdjlhlL0YrFfuSBkWGWf6VBIV2Z8b1XFCDu+YtTcXGR/VhJRT9xtZHou8eaFs9q
zrlQo3n9KrYfsOOl4+OAJgwm3N1ef2V1Cy3ZoncUrIDsmUk1JBaY3sgchqPJUNES8uXnHxe0fHzA
Ytcp9NsZdJ4Hr7grlQFlFMfb1Z6sVDebIUu30HCTDUj37e5BW/JcqEtLO6qq6i5KNUKiuF7Sjyvc
JjIUd89bepCHUT6eCnrJaEGbYnUKzgIHgpb8C7m31BUeE+NG/0cjMIsQjA7hrdWxTC20NKzstwZT
NRJBT/20QC+70+BMsUnL8dZ80//tjiUdOy7Xr4QCYoopDBUyGDRHeiM7NUVPnmat1HganmQGv4vg
xgkxPIUo4R5U4chfNkZz99ONPpKZ6tVxckkCDuTJ/Btv+VNwSGLTx36S3kPxDE2ZdCi5KDX0h0oD
3MLuXLgwEnGCqJAiYnUWh6NHSiCvws0tvR3zhDmZWMbWxefIR3t556mNKn/PyPxkvpOMVRFVXnBh
RX2A4izJs1uYtBRh87eeVhRCvscRMdXWg0Bk3mupRwQOHjOBBNcjjRwiuR2viQKl6yQ7Hv1BbZht
T8WlTx9XV9tjs4zgYngdSW5duLLPBhIf9Ceaf+dbZd81gE1CJM0dn5P4S5/16bG9TRyIRXf6OcaY
ds9/xt67FU1JPpnWJr8vF8p/i/ta6z64qgwUtjfPBti2TyLRYDPmo17cNBSMNoW/GIviqwTG2r0m
L6UdI2D6d6e5z/72fzsQ2Mjzv3AdFB4OFhTgTlGrAPSx/SZ2I1Ehqn3iJjrePxcHrTET97fQOXfv
2a8CnyNiJWFPxeGvaEVha6loiD94KV0LQQVuQBWfeGu3eyNgHRwxv64grJThbjPdWGiNY7WC16T2
68VvXnVBgJajJTVlQKp0hFGm/lInlB/qIHaznaIhNVj7r/RD+zjOP+hhej56PsYREhDjKKWsRo7/
Dsllh9FDAfA7kBNcR71fJAujgzm9d6BCs7VzDiDAkv+3I4Jas2GrcxYLrMUofS7ZNyhaimmfbTjX
GES6ua2Lp2DNnByjSB0aSLEstnhki0C/gtrX8VznCoGo9TSjCRVhBCoPRr303Ze93zE2ULFJp9TX
T5vhD4Uish7m+KCaMft7yRCuDEQvLYVlWpifgd3TMD0++onFGGQFWi09IdM2rznYC/6kWyvEDeHN
Ki9z+h6Y7Rvp80v0Zq0QEdIoPTqpnidLC5bz1vPFxcuLLenYBeYX+4JkvvK1/5Jic9riTWcFA2xo
Mt+9ktLgJc2KWpG8vP3ODeW/q95Jw3Jhwj6Q7YZWTOqwv2NMbp6EpQgLvQmPdQsVMGW+mQM+4eN3
rg22jqhlFKaAFvY/Xi3veVCbonegt9qWvFXSgQbA5ZRLLr9PcRAVam7vviGx4lxoh5bl/9I8TVjc
vA/IciWIddAWzRQJ9KOrxN422aX0JE3QUHzaLXKnxFtJCbazphzVaDhcgw0wWOTboeND6K2Ap74D
cg+ruYr8FlvGqTv8TLWNBlFylcP93biydoObnuYxtG6gsMSOwlCwW6Thh2mhiUoRF+VO95GOTR6J
PMSlLvk7ysyvKSjWhWGdKzUlRiyWbJ4fQYFPKbU4z/Pz6jZi7tcn2PbJeVTzQdgjcInoaY8YiXo9
7eq6TPkKcCHqsGytB2Q+fjZ1TSkjwFBb5HqOF+eBHq4BKzqX8l/OHltxNzt0Er4re7U9oLbIAQwy
tikv9+R/Zg5TsQRxjqQpgQwar/HI25ZUWRs4/flfCL13jmEanW26YZ4TbiVoGOBB6OuwuqubzXxT
ZIJscUny7HTEe+1us0vHdTA6GPTCEPY1TcdOcY36ds/PYiscqHXvBdY5vK/AjBaN4LEHFOfokuDt
HOUlNNMiWjn6l2PajOCIIFOM+Gb0Y5qHNCspBFz7n0kLgDYyHwh/PuODAMeIvf//S8bPo8UZpT2/
r7XInjqVYRRbdqjx8THrFu45A40tLZR4/YeyiXRa3BYTcd+Pv6w9svnMpTtIAReq5CUAJaPrddRr
H9aNO4uge5KApybELur4g1A+8CWStp2dHiqCPJ22sVjnm1hDitWq3UwxAorhajZKBsGL+50BexiL
bEZQRjd+wvv6//RDZeu9z/l8PKLx3suRmcWm46TFn/22ZrKem1Fl8TU+4FDI05f6N+eM1yA1W/lP
3uwhGR1JRq21zAVW2Go54S1OYii3NH2jqBG9HPuJo/UwZM4gRpKcFX4FzFU/WGBIRsg5VnAyaopX
OgsaVIJ62QFdMi7pTFeXeJaE+DJ26MbzjPzphqxkwG389ZGSNohqajXgrsNJ/cb4j7ivFA1ywEmz
a2GjG9+KlHlp+QjrjZPE5jPVSg5cCdCWHyik0Y4aWjXRwoFktsfxgEZLm/ZiTzv1TvzVFgSGctpv
YXGDGTcyhxvVKCMOjVWQ/QXbY2j/ojDOYCK6VGa3EgwbgqhXy5A533/gA9tz6Mqz1I3G1RCD7Ckd
SYk7H9fZVAPH0dNE34TZgbloS0xRcu0ofDJ967/UFdT1EUP65rchNP/OZlit2xbLca93VCYdwm3k
OpK9dgDhKndIBimgTXEFgFk1mMv66+D8dw3iF5wgYm+3R4UJ7CSAbV9a66zNXP4qyBzKfKjA51/Y
aE+cWy7xBXqMGA3IbGUvqtFsnDHpFG9OrajoVkvzxFdfwifudvBZqu9R2X2P6zKTQLvDrbXVpqxj
4uPwGzY/9fHC3mUq5eQ1zBAVR2MyqIAt8Nosy8gvHaIgNcf0nN5oMOMBx64to7txIwpVWLiL+rfD
/FpXTIfKGyeNNXgymZphkZHxwCaE1Ps60Pb23vEKtl5PGxm0SSw6IusTR+jj8xCczxqkl4JleFop
vYnSgzQb4mrhW1uiQK1VS+N2dQXFh7DeCjenuEkr1YIcaMz/8ixMoiYI2sbdgLtVcYw4zw9aWMz6
EOXBhJV7D7Cxh5s3k5iKj3zlc2TZEPO3ucd1Oj6u7u63lcllgf+QPJaXtYtbIG2yhUTWRQpcftP/
i8zke/JwzIyexO9m8udQ1wa6USYqzMT/YKfMDXsH5sGDN294mmaouVKOXslkQ8gdtQCk94+zV+DI
oXacBVZbw5BdxDW4yyMczi6rELRXehoR/Lo7ay3eZ+RE74T9p/FIZXDgiNSi7I0azXYybVCw+L2T
b6LtKQWloksR2069YXQqgJojukN/KUdpUP0y2dHV++HGbVDCMLbwV3Kbc+4ZawQjyo8SadQk/zKw
aWoER9tiHfoiOmlOhy57BFfcWeETde1zvf1TDIGdtHxTrH/i48YMj7WCsBecUMtxZcITzGX/oqbl
OFHCt0Z5oLtIKHFWEFrHM8UCKG3u7agv9mZL5sUe0O9jw0WxZ8+GrtU47B8+ZVpyLkP/u2Dzbkh5
8YCn61Ex4e+pNpyvogKx7RccmwlUvQGwsY7kZj6qd7h/A//DtIMjWkRAGynAFSrY5gw8CCpyk402
x2xrf01JFgaHRtBeUHMnjL0/fASnByaP5H6VrytfsKsHL2vAOCJ2ePzuA+p+3UgnAR29xzo7zf9R
fDKtDE5A6D12st0ACXg8fkFPbX8UEs5SEgFur9ybf9Bld4VJDCoz+JQfue9KrOqgT51rad7f+kS1
bQW0O0CxhgGDK3H9/adOvQpqnh7QlNCtPm1KS68OE7pyk+unvCUPKrFFJei+hH5wj+E0uLteaqbZ
xGIvj7mJlKDGS8qTExsAbCu70FZ1kcYjW/zX2uZQ+IilgQmeshMc94HlYLhTnzoFMNcntIHTzYUv
UuivER1BN/2NN/d5x+QzO4fW+ff5DZ0np+kKQrLksVMUROsjNOPXQgZZV509uMas7N7MLE60D1A4
bF1ZyNtk+ZMxc//+Z/lkgqcW7OMQTmSHjKQqMQsfdMq4G2w5lp8zYeX3BROz6n2C50+NacVuhLSE
Uz6pm9iZDMVB639ZnHAiSE7N0DVQTBNie4Sp4b1NARDoVpl0BPEb0e4FHJhMPnFVgISjXQBzl3gi
IUJfvmKfdbsakqci0e5/BR5HGGDQxkLCGiyqjbpd9Woz2w4XtedZOJUWKrxiCa3rMY+x6VRx4tFG
SHHprlc+m6gw1smF9VhP3fWTle6/LiLTlzC23a8lryOZtz98JMd5+xdP4UTiWOsnLl5MKLp2y64c
TDLjQ6iWJW4WfvzWztKV8podEofTbI9kd/jyUMgvVw9Xx+XWAbgYV/rjVtv8envJtTq8a9Cla8Vi
QVWSIDFhkEp2yXkku2JiOuCvugw4fQcw4NCeuST7F2dvOglAYHVu69P5iWgPArP15w758DyaJddA
keqIKpnk696Oul0ZcnNDLRMEDDnQb1AN/6+MPV8nW1hrED2gFWdFeZCt7dEDb//pSD/sKe/2PWij
nqW10itFNxi0cXuLqgGnqPIB/bXARBEh6pWn+4CJGm2mRT/lc2aG6Tvc5NP6sTliKGVC7lxj4fu8
0/ZzdMtJuu/bRM0A/opkdIM93IIUdvp67eCLeoaPBtgS3e8exk4WmMIzWT5+chPRcLqFTjKVEpX9
W4Xup6wNdSM5coUS2rnBWJkxzvUF/tIaEdiQncHqXF2MYVEPmkcZ8Xcl6wGcmF0bjxE4M/g1ryJo
0INRCFL8xS7xZSZVX70vwES9kBI93BFnmo8Sq/xHhiqFVpGb2gDvUPqN33bTNwOrpxMhIGCr06WN
1Hqre8QcIQ84oqQ/voouAtPi5PeKWrmEME4Eo3wluMFgqA9qUiZIzLoquOm1Z/2T415gEStqlH1X
J+dpg3mQ2qAftwQua+agQ11tGB9xJSWsjOgvGxZI2xLEf9mA7rlwDyExBlsDVrRhN+VaSOWUjNQ8
8r8MFlaBQ3rrywPbfMJAHzLQg4RjbNCQuc4g6/4VwI/3w4nNSIICXADDVf1uVYGUW2IG5n2ztEkK
NH+G23G7y/cQBVL12AqHSWIXwISgeHYopUGB3aZuDdsM71B1CAbMJMZARHTAZ28md9C3IPYXuQ2X
l9pMV+aDyebJQbmrq2TKVbY/6xJkOiy8cbTBm4nkkgXqCMawdyklZKhkSWbb4LgKbp5DCcLjxXcx
PBA0Btj+4L239WlIbtk58faScSWi1KRAj9q7/a9VahBGLuPvEtDEisaVSmHbzOPrvSld1Q3z/mT8
VjTzkNP7bk5ZQqi3lZy8QEkEklNDd8h8dhvDCBx1jY8BAsUozLyidu5fW/stLoZRFHQ5+aDe9Mm7
sAScgGhrd8PS7I4TWka2bdhHcjeK90DWLhQaz/r0rzanUcg618g2+JWJrdwrAUaXNjjFmsmsAuTV
fTZiC42xeEDBrV5WSweaHcTlSdsw3sD8kvXlJxg1h+UPTZMTLeax6zybqKoWQG2VimBWwPDh0/1s
Ev/rAE2p2+mxzqdq9PzLVidcf+tzluJLGbnc8AJEJQeMpFpdlaC9azA+UKo9ODzDRrChHP1XbAv8
ys27TBiGiKGxmF7RU88/AKqyNOXtv3/IYMfotmcQVzJl7qZbD3Y3buuqqEnkTTt9m0Zl2exA3mjz
UAXiI9yBepE6NVev7GehWpAGP0494leERaDrSRLyeCPgyR8g1chG8P9BPh632QjJUiUhrx3YuQi6
UBN8fjf6zYq8mkqaCGPQF1JpbteYjAl/USAvCWK2aVypFYskmahMDki7Asjmkm/OHSf0D/cuGsLv
r1T1VzTgU+tTnGmVsDVd9sdF87I6dq529Z1JOIS3Nd7TB8wKpHAAsOHnYKW1e2TL/TerwU1Ac0Sk
Tux81MITCpoz2VAT6ogSkNWkq9lZ7CRfJOCjl15h+DEhqpfc+E/Z/EwRg+QOqDeZ8JpzEuhF+nOy
nmnysz5hqMPyTgwb+kEufB99XwaPPVgIDQYt47sxdnKLCpAeowN2qdtCIIKIP5iokjkv8EnpTpRw
/URos40xjb9JyOu4TgK2usHix77jgwDLjWILD8nFwCy7pmtPh0QXr3U7rm04aE34a46q+SycHlnR
/uG2gGP+boTzUFu/kralIWLbJlkS39pBThZMvMvIcJJO11G6a24RaVABFlOi3m9CwwpYLk42vJp9
vcBoB1Hf9mCZ9itp29V+TN6SHv5pB4zJCdqiOtykWKVNBRoGYsXlS09URpJpeJwXbfkm9v4NKFR3
4qcy3ppD7WqRbzdDw17iesz413EK6IPVqWMFbgtssRpRjsdlXjWtWv8kfkxLzVr0y747vNM7pVGa
QCU/B6BGkY0Ykt0pSH3IJyrJMK81PXuBMZhlbv8kSuMghwlyTi6rZr+/ZOkbW63jG9BhW9aZ5IG4
Ggk8Z577ueUkkUSGpCzxFGtMisnowaEgVoyF25uaYQSAAjlIGRyGMkWbSXtHiCAVImRJbexuZQor
c6BuJ+aDFSodpLXf0tY8FrpwaUmOHOwEe+uunPRpoC1vwmZwpRJHShmHZu/vGrHJZwc8bY99MrVE
UblpXSDbyTZX/CKF+VPRSJe/a4qqkGW2dOy6qJ4hZT7UTMF8Hv/+WfXe4J9kqlEj0adRSKAsRRYk
HNxAYaBlhpe3LjsYmpUN4AtP6YuD+ZRiOCGX9AA5nzlQRJrFW+ywd63e1RxITElQzaT/iWoJ+eAa
2PKsjej8kGEQ5QfVUM/auo+AMt6LFLtgoDPzak9oNyaDo2Q5iH875DakKG5yygNAU6rvEVnOcF8y
Xhrv8weAmHdLTMZoS7a20TRLdDXhek4LshtttwD2ZjpJJ9WZ3Z6bsif37RhcktBcMzICaD7pQckS
cQI80hyxewnZKoBsgKuJ8YYqX903yaqfLUn1+phCtS3Z+XTUiAEXkVdmu8/VIDQ7uvaSOEihQs4X
T2/r6ufH6U6727qa6kmzLo2NpCmkxR6hlje6uM3wUjjLmEWHuJykUe+yws3qCgru4tguOPyV6hCb
wMVIJKNkDSVgpXubox+RjLVqOP6tf3Op3QLnWuKa327uhFqFDllTd3XYw9t3Tr7Pjnus/GDeHa0o
RlDWVYSMq2xy4c631F3SD+efCrkT5xidPOCerJLXdu74vxm2MnR6DLBzYS/RYGXfnfhqpKeiBQF0
OSstElIr8BQKrrlBXNsuhQMG9lTJSri7HI2+aecCRgxdCRG3NAiPkhcWm9+xCshsqj1xPOkdvMeq
bonXLid42vAu+TVbxGU8mTBxkUup8pESZwOJeMmP710V3njzecc/EIn3jjsmegJTGIDUOcKk8RA2
qrXn/sF+yXLCbniShyk16nwfLXpoKbGu7RCJ9nECh5/uOT+0HOpi6uyaf4+vVmF894dOs4diuk8w
HP1VHBLbcizSxm64qLgntCV/mLr9+pPSzyc5MOB1UqNqGBpJ4csEMDUSsg7MWYeJrh+/V8LA7hNc
c1X5nTRoDFv4c43tufqWXozoxjLPJTDTD99w0AR5ctPQiqrKV7badMmzbLut1qwHj/Eyox3FIxLS
w1nM5NyVLTJInVzq3Dfyl/EFjg9eEWVO1ssHFJRc6p7kzOzqxG7KOmWUC7lKC+OYtEarxEga1b35
sct5EmlftWvLg2khPs5XkUFs8eWBgYXGpWB27yoU+zOpXXzAkjyTR3dZ2YTYpzwpi3t2w8aZ747z
sLUopoouIEAgt+XxBAQD9nJBNG4qqlmvnKOzNEkhbnMoDol+G8yWFEHJaqa+O6/Tn26gFBVpTV+s
Ovm/FYNANmIN0SKsMAABvuMyM/nKEE7R/KHI1OtiI3M6AUWJibCSXN21NQEIR+vNMyN+RE7AuaTM
TqMRSnAOxg8aDJfohvFhQ66DMbc0ZBYk5H2VN75H/QfLmORa0H12/8vIZZgkCweBjxMWya69XKf3
bUEPso/c5etr/ifzBSpchgZ/8WyicAYme4zkyT0HNXevwJpfsqQ7op4tJ3WRizaWEdmfno328CyF
rICUQjmTcfzMUcRyaecQXJD8EPKv+dZ7WQGU3o9aDfkNo3+JTuD/JVPV83wmLHfdG7abunRpmx1I
s3lmSbP2S3xpbV6GY+d0vEO9srVgBth66oSiH1lyo0sNhqAY80+IYO2gcXCRAerbEPthOfnsyzQu
BDFTsA0Z++Iz7SK//FM8V76t25vHoe8X275kzr4Jw18vQCYrLPYdT5yWmeCld6VVdY35q4xAPS2F
H8jaY0XYbaM1oc+mm3841asXWIH7IV034S2gnwmUE06xSqRro3nX8IDDTsuYK8uB81AkoA+Rgs3u
yg9bp+kIFb1Z5EQyRwPvOXVslSlxpJugtIGRftlOpYIvqva1ZIZ2iTZ8NkWaP0R7iTmz+xfPMxV2
oo9YFyKvay9ERrHul9o4snI2pjw+Ux0urR6D6hLyDDhv7tzPXbTzDcrQ+c9XEsv7w/1uflMdJxXk
f0mk2m0nj8GRHilljbPEi2jk6qWf82PuUGPpsQlhBtbGl2NnLRdK2at51m3QOCNltLzrXVlwayt/
qPznne/XAprzMgfSwuIgj44PGXp6yl+AUmCUpPyqhEzxNiG9g6gphLOlt5oVN0iR/uOxkCoFxRU1
AxT+8xOfcdyYtvDUTpgVM2hL3D1KVX1v1Wr+hXK3qZI2x3XRlFmbZJcKsXrtwRLa9cawv50ZYzOn
zSyGgDxhT06/1Kk/apnO4Nal+0f6oKO/HDWGU7bNrQFN40DV2dNtoC5lSZ8yhskVF1WJbQ4TLnfx
eAcRdcLUddSuxoRxlmmpZfAlUdgAKaPHFWhRU66rk6Z3BHA01Hdvi9HLl418YhLYaMor3nP5PfpN
ZBO+OEg2WdNf+9mW1yVi/SJduzbj13EJKUhE7jJoqWSpbcWU+Li7M4UWJfUK/x8Q75A5mYnsWqiM
rvytgH3Uf3n66Tz+yZIsAGRjn08kL8ZkiCgmFFbY9AKtf51ZaKdbibpag7M+y4jS29MDL/0G1kpO
0CLJkOCivq51RCMxDFUx/j1s12QL20MI4vtjKGMvM4DxaZjRD2N6JR/LpgE33tbEPbPkzav0eo7p
PAF9lEMWOsT56n+V7c13EEmioYV5nv6roRNZJNkzDxauhgePeFzk1Kh0a9MHxVaRueEe+RKusvMe
SGFZulN5P+X5klpEr3R8uX5BJQzlI5Dmw8Lgx09+OEMwKdPNirvT+O/cGWUb0pPU242MF7gAQzJ+
aJzGM96vGErxjpeA3wR516KJ4rlXx0ZgaDamNFSyGGsHkAMbCL0W1vaA+hrZdMRPh1zXCwmXPGQQ
dX6zwvvcKDh5wpS9ZDpyVJvP/OllQ5l0MfLv+fDq3bVnqj861wuFIimxuolorfbtiDgthrBdGhU0
WXgQPFLHjBcQWlG25mMPk1U3QE/GE64I73HxlvwrWIv6+u6lcRdhjoms2twQR5SR9XxVfPrQHq4/
7dX/bZgEjo4DbrjlpfD5XuulA9L69BSQLZUA/UHUrAM8w7fO/50Lm8EV6C61AJi+lelyIvcj0b3U
SADBlaijdjYyCFjnMQ+BSP+T8+R9iR7RjaGxsargsWE8Darqev1fXyMpbKU9DebLbR6LyURb1rjq
DZRMFS1bjE4mfEego5wLJq2J4E8+CdnjSKFvUQgMlxro2CAqSfd3WBlJdTiDKFwWKM64DFp3Kh41
4iI6xQZYPVKABRK+TbJU1mIQVkYAn0yG/fX5t1//OxiFloI2MN+qblVxl6Z2X0FVJserJQCslhIT
puQ4O8XgF25Ksca/e3qUl1ly63qYQ+F+jyStyOC2HuT1n65EV6OGalFqxRNfoxyzkqQ9u9+sWsDb
BuXrVPy9qzHC8WbIhLBrUCVOFBEdVC7c/0skdCzR8MktwKNjMQssIg42b3Z7hNSRmi/HK7ZP2jr/
DR91v05ft26deXqkCDWfwo5SGBnsp1Pvt7DBzL52l9PSImWB6cg09J+Pu0TmIB9bFJqCCexNEdPG
giu+E4VnTZFeP7NztYu5W82VGCfLyHipw73u0hZrZdeySl2drFFuKgnZH6n5cmQfHuyrCIQVG6Oj
zrMiVutTTMlECB2blEgmLgoNeKLiR3px2v+WZEqtU7QT0wY9EySD285Nq4RtxATJoXdoMMJS54Ca
2puKQqrRMfwVmJNhbp6goeNClkyVtReU9iWHrgyxsY016XswxKHTDeJ+KWmXDxBBwhonxK6LCfG9
uGnkqNEmHp1+qFmE0+pZBLTDv6bFdjhnEIjftI+iKNvJbgVMZLMkO3HFF+i0baIyjcOGsH6AgE3G
57ILCA4E419cM/wW4c5mNnhCSQ3GQmtP7uWO2qi3ZtTxf1/MoSDPwCTKs/0g2LAqAkE7tK/lKreb
indc0388QNCxKIR/7mxbRN82wB8BQPIMYHgXqDlvfV4Gt4Xm9tTk/ghM0nPzr0QA5VQlnrd/4dZ4
mAM4J4+BJk0kPZhtbWyurgwg6dzK3M/6J8xQT59oF7i6jgyHClulvLmoXy9/H1XR5Gm67NYYeOaA
KhqEAe4g7D8wAXaV5TU8SXoN6p4vVCki5j4/kBjgP1d+E5jVJZFAJqItykVAIWHh4gpGJJRnOFvl
oWWncKFddm0geGno2C2LX2v7xkSn/aeYQzCG/VnY/FM4oDL/9V8Io0cYaYgWKXnM6Viz/eIvQUhR
ryuyi7c7iGvAeOjUCbrPfZdbWYqgw2AQqo0nXtXAgLiBr3W9iXZRurIEt5Y+uDhvnuFJwt2ph4Xh
OjkP+Yxv+KzgEgaVNGgTVvH/uw5pc+OE2Lo1ZDOUvPjyojTfSpi4z7ICzGVp2kr1bXCpe3wEQ8YE
9nynh1X8n2uT84NyydN2tx+UWjhxIKOaEEZYSd2bdhVOaiaSej09pq3lhBOBlDUZSTla5dUigDfX
jQiKDf1QrjuJyNtLkntDt9v1Bge9SqfRvw0Yo4CHqWvrpeStWGdcOgtyVOQlpleHcmdS+KOxAkO1
GSGCVTHoOGkWpv0KPq9/M1ERE3SgYv+5JpzYYrm7BC3xk7jyKKxkZ26neQg5LWQvj7iTaqUaN5iM
8yf0GCdgQO6sAOK5bEsNG4RxyMaXH3poWXLT1RrX5HTopzA33nI2o2veMYSSfLJpGDVYeQgBC+Ai
JpKR2+fyfitTKKo+bL4sxKTHzXoUtTRW8yqdBPsxiNRZyDGEDYXekgbNsOIXcAPY5ubIopZCRuea
iJ0DQMJda9bllrMJPOyNArvNKGMFfbgQDRstld0Cr7oXQlfPIXzIeZQJ2jy0sToPH9Gqb7jEDL82
F22HZapUrTZLmBv5cBNM9hke4U8JrMCz4cPQK99hS8Vdzk+14PGToOjkawNinvQJwCrTbDAjYV1d
KMGyxlfX0AYvOlAMfmq3BFh4XD3PNXCFQ7VxYvGv6UZC1mBTn48KP6DFx/ZLCaKiaEHtjMPcJ91W
cvcifqwOuO6saEqzKxOgQRLJvU4+YN92eRJ/gtzh6MNLvCf5iDnniNH06n98qnF5+yoaU1ctxIqa
uN1zyIBlbSkVe9VBzN0qAHtlx5xhPzwRmXYC4ah895++3elx9CCG8K22u2L1cDGZ9xI78NSJot9D
JMuDF3A8yM7JCzANGBVOmsGRmPGnJ+QwGtgOq5jy2GrvCCMe62R93vRxAoVodTSuHpV/lIF4HN9T
Gbz66x0Q32qjVjwGcK3qADKv7LfpuKXcS04Lcsodb0ZqRaxFoNuWKx1FXzRwDQiK6a8xRP1uuQ2V
MiXEmXwSNSbi1X4macQpQ8uDjMliXS4Khs/LmjH3F8h9eng11jZq2rIRfNmJR30x9yYJxGqA9qaX
tEnEWbC5lUawfa+Yt2JZev277CmNO08cADVffhyVy+PrsFj9Z85v0AAQqTuu+GKQKTe1C0HfviGW
srE1pe58OokxKrKzhN55IDYkpOObUJzbhDtbYjNWpmCtGGjRf7pGnXFSDkxGIIHxtcJyk/260bEC
O4ylsxMuZjVB5uEFl5wefSIDuM51zNvgsXcGw2SLwHM6UtlWLHWvXQ9W8BafrwGdZqTISgXiNSlV
EdUdWjfmafegYRsjdZe8LcCWj8R3w8e4TUDpmX1rXDiA3YMSZx5Ep2PPW3XDoHBD5K5EViB+l3lM
vAqO+xcMqmzr6PGJ+UgMhYNNykm63KoJULIXkEF7UtDj8wg8H3kdfUlpTPpcybgd+MpCNkFuPEbe
19xUTeegKPiEq+QTkRP5awHLG/QJitQk/2NyTcHy3GwxeU3uTaQtx+Q9JUunZzFa+DmxwwdshhPc
udp1aFcvsRDUeDLqVQto/pWqOg1CN/XVfQuxoJGmv2qruAlP2ZgK6jxfeHm84zjGVRPl3yM/626K
qAY//27+hLeVz1ZHtrb98vJqN9cMpNEZASa/yo3hUFKwHMWxQwbAACeETH2DzW7p3AIWdjHlaUf8
Drh2TezcZfs4oHt3f/SBLHcLb8H0FQlAJntQSbft8SfwPTlAzuO88c7YLwjX0+hmgGKIwUxp0itW
g3rHZIMvtHdBorXHxjd+XnoWm6u50t3ULBVsGrRbQ6TX5J83w6rMf9ls86kUkd5PCFPU3p7Y0k/9
AHbuLLsit7zNjWC2jM0NTtHE7MFAYCninWyjdLanA+eJoX7YH8Woq+DHHtexyMYCRdZjZH5syfBR
4dWL4+80FORV6m36cA0LkbOpSBXuasYuY3khb8Qz3R4LMDKMZ9N797S/MqTEOqNwYylzAkfB0JRy
EuB0zd3cOnpcSaDediTLgUwR0ncfBsKYmofAphdwHJzTWRnnKcfFv1ncEbBzKpo1QOzyPb+U1Qeq
KyX9JYqT3SAD85uLElYyAc13ukp1H/5iQjIXKhmchxtHrBhyEx/6RHaKDdXYP1cdOw98TYcS7y/X
xs9lbTrHySI3A19BkSCDcMs2se6BZnkyHKhsU1gu0yqqcezmXPDa6DTOc6ORSbLBL+xq9ynu8lUY
zw4Or4reLYH8YyhcVxnkCr8QDooxsZzOeeM33QDCjpfxBo64WYUZtPwVhigI/nZNZWNd1tJH9i20
ufdNs/bwWhRNOCbNBtpBfdadDEnG7Kcava/BZZsn5wxnV1+hV14rbjxt3QxLpqXYuaDvPRnYliZ1
sQ+R5tFaSWrqvou4Q/4Y2IUdpdqUl862N+rOTxSTni8OIjH7AyO8TuJHzC6KBV600EOilEenzD6/
NYEaR8eQSOrKcl3o7f7ebAnZ5MxispzgORuDtPr1WnJRcY88Jt2CDhTR5ZJXxndgLZ2Wc5Xd7Jcp
vzzGvw38EbZwTlOWsCxH06bo13vUfFdyMWlCw5vEdPg/C7SjJaAjj5h+jmv4bGa2EDsaamICBgVC
k98LI+sacty063FD9U93FAssR94jVdB/mvV/AWM8OwO7Efq6tGdkOQsP9ZXG/rIY4qbtEVBMIsV4
EksWmpGWeD0QbpAQFpWrzfr0cz+ajINsy2IFGVqIOCALo/00dWsxlFIxWm06RClJ5RnfsYKFHW5u
arDuGZfG7lxxfIU5eJ8E3i9SJfdsguBnIohgpIiTwa/TrtgY+tb7cERVuvAfB2SjIrLtw778/1j2
BCCO+bTLbQXKudDECWYAbi8fD2ppHcwS4Eubz/r4NGZs9dl0C7CKmFOrh3fVdlCs97hxJTiOxE6K
wBQXPrViDBK1YxtHCEs8vxNDJ9GQgIu8ai6QzhSOHeCdw1cPPxnf2ai9sZAO8VadEM/24eZYdVNU
JF1kwN5QOmuLAojhubu3sm0Lksy+GbSEoD9NoJfDfKytdMivl6+kMt0CMfkztaJGvJB6Gb8J4U/q
/DPQOQasjbl43t6q9M2S3ZpEAQ9hh0MzL6vn4uOpC8ym+sEFmJ73Sz9rWVU41vA4OWMvAPFx0OOP
jQiAkGTDflrT5gufEAf91ryg65N78KPq6DV5j0XonpfedDAtLGTlW/lbSQFBpRUMgZzTIfJ0XrnT
t94jkPdoKT+FPLr/E8FtkUofZrjmZkbeLICeii75DeWj2no/gQw9LOUt9RDN1eC31CjjzOpbXUib
qJNMeNdaKCCZsZKP6LrcuqTpDta4aXym9/YEN/G5EdN3QJgfd4e0F1tSZqWvQ76uNp+DKgT5DKKn
39w5y8Z8XWZoSXR99FnirYugxb0KOxyjBMhB2MjDq2WHF7xALSR+oujSgDRjNxrtuyslNOVkqHUo
I8VphgjPJgusE2tKhukI/bjBf8Taf8L1wo+DkUOHR0FMAiuoJHSJqU7sJv3KRPnQbSICwJRIApH2
gF1D9mZRkyTvFZjWBTTXIFufLYX6BWYDv/WRN4y/cpiX1+lFsaN+kKGWJYgDdMfU3BhsHK37dOAn
LK5FJm3RhADD7RyYnWMFoopLpabJk9QOGvbgLUIuzZWQr2WCNFKY+Abtt0mUXdhy2NBmUYvY5qw6
QxMqPSn7DJAdUe4MWsJVXR+dGXcoXujOZthVyI31mzw/ewsuju+nowUjXSFhrqO6SyTIS8wC9Dyx
85QGHkROLTeH/y0Yt2GAyiyNudPGtM2zIoUgddl3oy5tsKp8m/kar5+SEA/1LTMEWfWlG/qPbqBu
l0tWs42q1ZO1g9IEzzVqZR2h1ZaLLZcpPC/Bozw1Etn11b9Q2lcpvdGVlr5/DKwvIa1jEt2fxPmU
sxwCun/7t7+LAdo5bP17u79aWtiNMw0BjnIEua5AQfvkgMGXjGLzy77NFpARPwocXpe7peqC8e12
Bo2KhtujghpVI76uCJxYjmW98F37muNA9vrTwPqx4+3k+wzxY+pmsQ9xf2y4OaZqQ7FUaKri7JyS
3ZWSI2SGffQKVqRR8bKhjr4VN0bhFuNBmxrQeN2CzpEccA7RNpY29sO6qn8QZKKJW7cOOhkcrKwW
lbiqqfa9BkyV5G8DLbMe/AWRVI6Qg+U0CCP0OPuCo+dEQHPfrQe0CNFhxS0hvieB9kGzyA9GdyDv
4xOp7GnJzKvK4tfW0ZebHL8bS8fKMqcHNUfIe27npl8d6cGOM4Y9w5elmDPTDwxNfgFHwTSupBvv
1dkWHHiZNEmSElNnFc1pONuwqpk0XxE+m1DKhinIadIz4KjI3Gl8SYYSrn0oKU3xk1vJm9sc0IyR
eK4PcqDxdq9SUpUgLguA1lbkjT2oQreNFRZYf5Z3owSLfHp2+Lm6pfj+3HGTVfou3wYJh9Flc65r
gzC84B6wlidGEUgdy1r7d0MomscNMj0jzrbMGD13Xnh37m5c+qML9VUxEIoskNgz8OG20P2IKFZS
/J2bgVBHpJxiO6w5XD7+LvgboIG5jRSJoTnlg+oQCI7teZNAYQZtfiLM224nJUg5U18y8Uo84jQw
FpMd1EeRpWqwYINZYhdpOe8Jb23dH8DwjtA1FfjxKWISY/Tx6jA08luYgRYA77eHmMbz69kOkREe
E27sewcVcijuQAN2AHARk8mjzAJnbbM03lgdgPN1y4xWe3LDXWHdM7ALLwCfhNAX54h1R5nRhss/
cHPMOozVQ5ZKdkAULyWsCkoZ3cZDDUeB+l94VLU+PWfrQKzYAgMzfkgdlc+838MN+b1FybNDkmNk
UgkoL3q0Rv/jJw4nzC/bp3BQLsJqjkqaIrwG6N++WNkCU5YjgHHBQ5nmn+Y+ZGRedHL+nEjVM+Gs
fGQ45SDMP8PQaqCElN55KKeEcpJ8ZKySTpEHMPyDl0SwxWzkHfcvncjYlWaRMzHOpxyzFYrrb+s1
mElSCR5bIRu10+1rXiLU1Zj1ClLSdK4MeMJ4Wapvrn27XYvSz5S2DlDA1ujI0tOViMgu5khL1zz1
pG21ZsaDz+z8G6+h1EJj/dw3IhxFjQD1N/KgA2Z7lxQrgyTA3bBnn1v5u7dD9NczQWmWw11ChsO8
4y9lFaAmpghnIC5uYwH9FCYgGspMfNPc6EMKex2c0WTuj5eA2WClZffqw1ygELPaGAGhbb3XApwE
xSYokhccR/GXBKsMByE3gWB2htcSyktUv+Ycv/6Wrc3GQV/YGRcobXSikYqvXgWswV8ZUWtJxCbr
FZXqNl3wGKFMnQHOzgglScj5mjUjmqnqO98XeSWtbnnjKS9u6iL2CmxskkywbQNlnILAg2VAMS9q
X714KiytZ1f46L7Ozhn6iQ/kh/i5HFGKKDU8X+bu36v2NxXtua5YLZK+/+IidqvEJVcBX0JYVv57
BaXjyvkczXg/SJomcL7tgXrVrRt+vEC8XezHGOjd86dZmz1y8VbxcjeWze653L0/CkGwR52guWZJ
7QoEBHJCcYKX72VPl7XlGY6J8ilvWUTm//AMRRRaH7XF1kq2hD4YoBWbsmA915LcCJ3i93VfBlyr
HOcJlftQfjmpwqlzkFEfCjIHeLjInAhLndXk4GyoSmwcMw305fFd4AMjomKq3Pdxc5xy6mavqQSR
p8Ezto9jMa0ZzhdJVe6vtOjXxJuk6ef7w38XxM2NFKWSsJ1NOGym8Gt/dZmCEjF9I5gsl9iI/xw+
7RBJTy1QtVeACz3huYpjOORvzdiOzffWPiDxNwus2y6ZJJujo0EVdPnBVXcz/gW0flRp4zStSwWs
9eXMP0koKZFyNcCYwvaWYlu7hC38BEIXmc2r3KU5DeBSQC8x5ieJXzvKJWSd/SEYcCmd81e/98Wl
J54crRBVA72feGJfa/nbXzu4XvnL5n2LOWqT0r9kATU4MUNCjed7wb2vBb7smwBAcyjCKJW23BM4
QyBpgbhkb+Px1dPPpmfI5QQ6KgFNWKtAJb797oq4qXqNoa+HW9CfraeODaPWl5r84LLi195eh3M1
KsYA1wOHNGFy5LJVoRO1WhIPRg8S8zFH1dMMqJadr+gU1yuMMBf5tl+T+92WLHf3G5DQbIZp697Q
2IBKhqAydfEpPAzoHtg4NHUOQDN0kvp2a8Cb1cgubv9Eam+GvpU7t5ACjSvmqIA8BBiB46ThLH+l
Y66IskrBKk11OBHowXJXfvK6ZKiD+gSvi3c6T1ICVHSuI/FsaKALa/EJapbwWDqiNwGGRZ11TqYq
nNNYBYxwGYpWQItqpAXalxyWTGOJpIqCLxvQebnTzi420Dy88puH3cz2oRFQFOkqDwEHZwcuerXq
mA3XEHF10s+KL+VXelZLeba8uZUXWo9K3Wy6eIZYrz+56hUFbufXq8QtmmCTOpgFKeXIqriRD9Uc
3DgE9EVXCLHTqlnIr5tfubjtE8wM9R10szqJVbTR/h3aYcaO5P2StnI4mt3HvGCR+Aqvx2Mx9uSy
DcFIAJlVULo7UWae49A4b4UJ6jNi0+GtL8ivEK/i8kEF/B5dVHviTCBJESF5n0QL/UoN9lHKKKDo
3LHOH2BOTgQ/rPGl3nC721XhclC8ZQiuiLO6JeDwjjXRxJU3/zD9xdDiBoY/LIbnBYyNSD9NaG1I
eOEshx8/7dm7KePAd4Mrh0kp0EgmrNc1gMOYE1673MPGAFPiuoVsJqnKvCsb+nFK5nV6AAm3PY4t
qBMeNsINFOZCvBLk5EjPHWPOwjfF4JPZd7xD/hLx6jR6D0u00Euzxjx5YvJMqMkhs/3zkLpSSLp1
YooEcbdscFCi0pEF8j7eKWO/+mRX8dNB2rAFUJjL1/Jk1NtIXztTvoPyH6qU/j0jULUNXy3o3/nJ
Pe6cnWbFuerx+0kCmHc1u2+3k0RTPsDDyhHFtPPLOJUzPVtgn7EPdDjJF6Qgh0ZujYrPsU638o0R
hpeuXQ0IMKYvDMeLly7UcYuDXrIJ4rENMHfnzNW0xxDsLF7ntUmwjp63qpWDADJerX8iisrsj1KN
GTCtkAWjtdnCbN5RyJzBN0/UXGHyQp9R3XaFfNpQcbiEtLcGjBy+3OV1V14BlYFJ6aQzBj3EIVIX
tTyIZRdNB7FTyYBrvuVjkO+rpWD0OLtqQ5E7j5WK6VfXutO3vwwgIwwaW5PkjBfThu8BUrIe9dOR
S9SiczhDRthUf2TaZdK7Ng2yY6TPaBf8YzmLLDqY221yxe5oPZmvV1VOuL3Ce9m9kuI/LSazK1B5
bgpq2zuiS39AG2ji5LbM+F7i1pXi7XDCQgYiZtfm1LVX23blIR4x+1gF0k6Vf8Vbeg3W4bZMUB/W
a1P1a9uEgv+SaUWBQzT6vKVtHLoZi6yccQhc0z2H6E9alG3Cxp/UgSuRfdqFYJ5RqMnbjsZ5LVU+
AhHdWzOfQr0hMjnz+UHrLp7OeZS7GQqxP3qEOIm5w1es1WMGhjhJf5X6Nl6Iu45BegrOJTt4XxMo
AF1a20sQkfei6uOREiLpZ389hHmofIvuK3apVoy2YotSP2jdaRxipjN4E2rIeN4DNMbD+wnUr53p
OwuaQRGczs4QBGlKuqSTs0QbftS4ITqIEswtXhjiKoSGGJXVd281GlPt+M5qBdH7nZTSAhoc+2ms
lclguPQfqh15QNSpt7ZO9dUl/6rHTt4QF7xvMNE5Pumz0uGMljpWcavhx42DxqcRJq3vg2/eEPum
Ww7lgs8zKSyEciWI0EGmiDAivi0KftanVuDdgW8ckxTDoNSJVAeFTTHiEYabYPm40YgDvN5TfNOM
Vm2mPuL+uz1++arKQeP7aK3p4TnSqBIqqjx2QD72CxFBqVhEjB4otK2c4hUOBfMpG1D3VhOjJn3o
dakOtiQBZ2ABZVjYhlgs2V9wwlLhQ/9njs50Gu6P0B8z+1MVCGIFwXuumQAeEfxzGbKJT3wN4Qi7
9aWjUkZgxnWScrp0wcD/LlJZkFigoK7Dp1zQCK/n5aWJTW8SlGhHo3QEbUUC/LnEaMrKrGBEPLEF
SZX8Zoe/xAXxME0KxQLLXL1QVkqG7EmY2AbpO9MKDlOTa+wmJWhcLgsQP/e0YK8NnL48CoEXFjd6
aOe6rzH4aZY8t2taRfvQltGWVpm4Ui8vPCX6jRQZDA8ONDw+//pzNbVZ6O+hLbwC6qF5ECj7UxsD
M/99QsA25YBvY+bCQ7ZFoNezxwCbaXCDDpoo6nBAQzDNUDRXANWU7cKfMQUNP8TRWCmwV0lh+8PL
219wCWPaOzJJC/NRuYSEgE2F1FCbDxgUqPEhqCcZnkK3VmAzcNj6tQ/ofljXSO8xTniNT3e6ccHM
W7omULyQKA9jeYLTb1D2QXjHLqN6sAWtv4ly0ClZXykPvF/Puj39u5mKtnC8DXbiCwCQ7NQ7/e1f
ecWwEsA/zAyClOarxCIyvgG3F1saIUPI2R77HFBzQre7f1H52aa6M8J3g9dDkfDIfawGZu0JpeGy
0N1OzHJovdrSaXidFrFSQMeUoYGGbJom6jS88skyTrOoZ7rqhEMH6o2kmR5AidWgANxji/gRxDRZ
Ozil3u08ZgEVxAb5oq/hEpcEEhF2qz+nGazXiITUKZXvwuND8zMHE4agne/YuHGJHW5e+kSw7oZa
huPRYIAjqVB6K5Q/Jnr8cQ0xdHDegr6qWfHhEcottAwZY5waTrHK7f1ucJKQZrLzoH33ZzR9VmeD
kcg7jjuL0OdpJdp4X5kjX+Ag/YR++SlJB09qb+uAkMqsxjHw6G8HTFAVBlR+Qe8cwaclghOWtFv5
GUEOxNtpH6jK/WExVHX1Auz3AxSu18rl4fa3TpeySbaLhSMnY3+O2UfqQ6ZVA7jxxSolEK9Cnjmw
3SkKv13E4CCj6u69p/98D49FVFAV/gMzfA2L9dpPALH5gx4nRixEiioXVyffxFLHel4MkT7r44BX
fMa/+Az5zOUOblUstVIheiFelM0lShOD/zvMI/4N3AM0HrqYljXwfaHs3fAZTD2bpmB6U+dZlBRD
//9HxAGkbLoNf4OqQMp0LT4n9w47/YPRrO3ghTNc+QjfJYqH4N9aDRYUSXm2vc0XKANLwqusqvIt
QPY664Qf+jhf/wUcJvuyaK/a10qcfG50J3ZHS4eWRTl/g+2KMRaGIse4dE1joNVKVgckHCDd+Ind
q42PhXDsOKhDA29jpEACUM+LbAR5x53dp/7Esos2TRHwuRfiXCg98QkvX/NTbePNjfmYZTSJoDBq
rqQM8obBdIpDtA3t3cCRT8ShaTi6cABKq0x0hOmz+4BwFvWf0+fE1CXRgwPxz1V1z2G//2tmdXl3
kF/IDm0f5WCfM964F1MFSEOYf/KEatlG/V0hDHTz7Z308b9TZV10MhFF/L1JQFyeRSojqZ+ALVCW
w1u1DdgJcTc2hQrBLGycGkXU7kqcvDTndg2e0ChXLN8ZEDDi2oYA8g/RDtGRCljr8M4MvFWuXvNR
yxbPdmUS4qoU3rRnTf7qlBrCWxUpSMyQs6egxu81p6AA/MgiKA2bon+45vixdaUNaMjBWF8PYLiW
Ssc8jc9tI0P2wOEmAbcNMDIM/liCvvlKREQMUIntew/VccZB0mj5lz/1+QaJnciUCm7LM1dJNOiG
IU4daB2HPENmFBwgAIAVmZJLAUDQDpNaKSSFMNkybBDJyUwzGUx4J9/zlqeZopROlHQX+MY94OH4
dc5rA/3HQe65kMj3DZgeTk+r8lxG+wcwdM9kd5J5bJ1qFXMLB12na5U2DapTr/xsu9VxonCx+0Oe
DJUea9BSRLsNn609KSqFwqRG1gU6Pe5XMJws0JQObApgOAvbFTNJf2RvB+4bWZUo3wvHIcAkwXDc
i3tLFRyPShH9eK+qtO0BQk148QJlU9i2hkG3ICZDguyplUTbfc9MaYHlz7YECp1GSiPCdxEJNVvd
SEKSmtrkNHli26+VespcJGgfgnbTbrKEJzY/CFnpgcWcrHMFSPtwEB8DiDaE8zfHBu0LXPH85QFa
8dD+w+dycMEEpxkLb9Pct5xVgsHsfgStjRL42Uw2+GGTOwdMqLCT++mmI+duh77FqspJIV/BXmBj
+hLgQ4paX/EwGHBndJl624Gw77XaYS05VzQfdskgpMj9yNdLp2O6OPQMJ5N3GoAk15OCDrsjzV7y
vDjKn6Ag2HXZLuYMQw/cArs3atiuIpJBye3bM2zxa1ZN7i30CNjr7C9h/NOaTWzTMPip6lm+eZjm
YmydXzxWX1+Vdl+aHoyg66EXkgvl55zeyOD1Jzfg5yImv6RA+LCMKJ0vNLqnMpRoNdJZoWVownvW
lj0zf0PWgfGYRAhhXvyr2rnu9MsaT7/TSpjvkT03AcD77CLWVq2mi14zaOc7vMdPXH6sa5Xzc8Up
nUSPWGIGjGN1p+wuzkpAWxPjLsGYbTak9+NL1MgwOuEz+bHT3sFi+RHAupt3zPO9lHAu3Lpvy/+2
qT6L34u6O+oXlhq1CUTbSySgnSzqco8ZdX9Kvr452o/Ebf/2n7arJxEh6gycuxvKd6bNd3Zxky4+
HfEcMJbZhi4Kpr55YjDGjwrZMd7DE6FIGijRyIgPsx6DnyapjBn7ZnFl/5D4uKSq1mgYeUi/r7eZ
duQYlO59l+vjWIu5FtDPzg5U5xV65awzNOBMxHKfdbJ/HNCZHhjH5Q24CeyGxv0wVpxt9+BLOlbS
GwbTOzWlOYisoNn5ZosB6LMEhzpwl9d7n2M9tsaTTYUC6y1+hsMSD2usqJ9z8KiF0ydprOjyhiHH
Ym3QWRqvDbKdUGGjRmlJ+2mNeM2Tnp1pfobqDwI92YYSy4YAYgHkeevR9QT4vvuFk3GN6nhp9gd9
OH+1IxesLaPv3XNSGLjvYB+Ug9dGFAvy37A6+LsqLg8Ldcs+X3TCk1oJxK49sIcEGHmIpUKqkuTt
1hTuoUY+XA1ReTUoBoKMAW0TxZUsOs9dw3svXIpDw0oJ3HPv6jhvDrxO/OspZ9gGEC6GPkIapbDl
3+ImVXFTd/pWC8j9UCIPeCt+O79B5ddb8pSJBAMAd76Y43K56R3/O+1Bn4X3G9ei5EFo5dVluByA
GkE+2LPZEHVTrywmgvhxrORP0Vvk9sMZ/vuPO0kLGk5Kmkg4qzi/+o1MqwyoDPcTnujxc2fdVB1c
rG1wf04X9zhoxhRZ6qcyZSpZLMGSvTbCmVRl8MwDJ59jy5J2jnLaEhKn0mUJApZAUs7VHzvfKMvL
412s06SPEwAnB9/fp841OpBGDPxapyVXey9D0oGHWmSO7caS96EMkyE3h9klCTLPPetRqcFpyV+g
gNEBxrYFqQucNn7lAEVzU/213NTi9hlZu0XJtxX0GtFuRpgRf4v/eK/XtlXwrZ/SDhzYWajhiQqC
ySBu17l2q/ZOmHTPlfNMerZRRoSRwQiFAYYsxce0rwZfshH7OYZXzmeVwT0eFNChfcY26Nyn3p2P
Uoa2kVOotISwDMEuSLqyDlefU5WhBaOEkK6XSQSEql78UFDEqaWIz24mN3B31hYhRyoXt7A0jEml
0fr0blCeRXyIwzW06zTO7XGrQM51TE0xzNt57aA/XwWMKxb/IBRb6FBFNKgk5VG/s5ieGNV3E65y
B69x0j4R5EEtMI9PS+hnID5N3J28L8tUzziONLqAApJe8YfV5J/0o/0EFWpDl+O88FtfHYa6WXbA
fLAkmJJHc3YARVR9QFZzfZKDAkcwvHN8cj4tQjFEUbw0XajAx/GGbvqq/gjI7arAM6vj9+9AZ7nY
JsnY4sP8AZCVgUHZ1TtV1ptYM7mPGeUgcE8HOnuhVpHQZnNs/twlsHiEP0urJjhQCE5Cd975czDq
pRGXMMMwEK3M73aPlzLSwhRFb418myFXI/G4S3bBAdY5hMNw4ByHsGTacI5mQFOLTIiEfFc/9xWA
2xE1y0tdTGqpSJp0GbM/KLMcci5nGojoolk6JDAdOxlLV9WV5yTyG56X/T7dBbd9L0LlO8nb88NY
a2ztCRFI2kgYvLGJBGXZ6sGtKiQGLghNt/ij7/YmiZ4EkWHz/tnzQwrVo0wca+uZUHEA2+Q2fsrp
ztjWU3C2L7docvD8EgikvmIuiUjE7l8km/oGOuyod/YrRbuAqaJSXxfTwWVQi1YuaTjofQOx0YVk
Mersw7w2I77kxwKC5EwFZ/DugfXywPYmUYEeTpLCgK9RCw+B9x1SrHgvK5ZoSU6VzVm22QHvirre
z6/sWlRYPBPlbGXvTmYClWNSPEfzRzOCZ5Gdo8pzAaJkNHwRUfLqCXk0XgoC0GZTiAas9LkhfQMX
d6R9pbZ4rdW17Jnu3XCt9iE6T2AuJbFtEb/961aN4+oksPkmJRiCbmlvX/ArwcQ2t3CtjXiN0NRu
Ue1JjYbRjZ5ZU4Pw5obUv/3P4tsM6OeQaHwqKJMaT0JIsunIy+t6+7fCJEGVV8zwzQiTRCAsOEz6
PAks/wSek/1TmoLDHr/KxiVyVgRUTgYZoBcPNEwZVNOVKf1TBKND/RC6K5PXlsn6v57jADpRdgN8
KNQ2kM76JZOwJlkohOj55rm8yC+w0H3lbzORlB+IpO2S7hQNjaGCrwN2AU97nDE0ojey0R3VkecU
xaJ9FOVTYZJM/gVugfApyQmS1UmCpr2CEuXDS+kqowFM4Js9xoDhX464pn80fj8+ZrBsWqWuylTP
F0229YqCOe31b9GJVGD6mHIwhuD0LWLAHen8rC3OFOYL2KJp8SnDgT4wvq5fRr3KU5zt27DkCb6z
JfLyG84HnRFCss2j9xNKaoZDve8Od3s24sVdLv1weWQ/JEQhEtu0BYY6CHrwQgY0P60GS98HtGU3
GLLk/1uI/mbXZyioQM7f4e9wRuAp5l0uPc3AHLNkye6bT4e3qPeLXv5wdiAfwgx5j9Xp5FBYGXE2
I6dKhlw8Ax7/s8U1HGHxu9DtFwvzNvt+Ro83mPC+X5yGxbL8DbYURaQlKec6hOuQibTZ4HJRaD1k
HUzDOadGHIZ4yc2yYXQi82P5OtvH9D4/73mbOMHC4TxB/tAcruxuahW6N77+trpu1Gzt4USTRwnB
HM1spELmw4/LwPMACwNqyl5ePeb9XtmYof06Q8CLRvLkDwDsSOX+pnUtr6qzF/93WdSHah3BjlnR
frXxeI3QAxNptCC9CAQevA+WNIzO8+dxW/rTwmbT5Xm5t0Zo+8286tomHYHvs2PCbNOTd8t+Q6uX
uEcpZ7+HjM2qam9ySbr6IyF+eUxIeJqpW3L34s1LbhbJLFt/HJHaUDadvAHZby1g1/vzqWoy5sWZ
bb8KMIW54H/7mNhSfcZIpsuMvHhkVg0J7Xa8SxRGH1WYKhpkns2OnnoQ+GSQrZJCyWNjFMfJPmTU
d2A443zBfVyRy5s1F3H3UsOHeC7EAqyoUk6TcRCUATUdnPHL2DDsdw45jGTYRjVtrd6yG6oebCWn
1x95kJS3r4YqCUNLa7MORNmERi+T4QApy0VBAVLKcW4fsV29dHNXCUKeRWdexycskTR6hvAhC9Hk
dxO3Cd4y6pcOvPTz6dHUy3LqAgPYKeg2Wo2DxhSJhurR8w/Sf8UXgS8LM3eTcTy1G/x+y/TRmtWL
3aCk3627pDRi3JGDOnhu6tsgteF6i8VaKRB7uA6mVz7q8qa7/MxMSG9Z86Nl1b7yPVr2vG24e0oM
gEVhtJ0KhCpwidzngreTPHKKGHLSRrYJPtht8Wi7e34UbC0L7dxWRu36QkskhHOOsH/f5+e1pAoc
Byz3UWIDF1HE3lGUn1JgVv9w+AUtcxCe2OwCHwmAY7yu+CdZnbPvE9K3ykstW1GVky9qIukcCC1F
hUrpyf9bdOhbSV7U9eLoEHDA4TBzVBQxT80wd81H0UrD9cutjVR/PRHe1xHOFeAYrf6HmLGx2eR2
fDdR+ul0Zn0DffV7gVi2UTCRM4dRcCMXoI6KD3hkqazM/SDgSZ7rhUC/KGYXhGjmq6tNlB3gPf1l
TIZW34m4ldyP12xptROcICKgPNuvJzzaZIp90iFAB9xJCxqQDsg4GxyfbpDhr9/ijDQAt02rfUWp
Cq+mHXuyMSJ1yyHHxYwC9UUlYIbaXQTdPYwXTg+znWrLj7VGIvmXsiAjVgVSLm/gLmch4CJFci1X
UagFe7DjRdFutD1Bp+a0ep1JCMT1LgN54uU9E44dKIsp3M3wFN821hNuquMwC50nl8D6sbU1Mg+0
yt9NqnVTKtPhdFgfR0+d/zxDBuqKJw/qpuRmZDCcHLKHGPTH/InLbMtpqHm/JB1tqknswnYsgWmm
2qSVPI7/hdcqf4gNysvf/a2Kw9HDRMXq36Id3rvLsUB0IjH5khqrbS1Kziwekua6zerZuXZctCt/
Q9BWPQBlT4x77Er2Ekg4AZZSJLAtET9Lvlf+Wg6hksrVUTJkkiStJ6yJV4ztWNIOggo9/sCrJcZN
SGvDrH3xeFN9PX3F6A/Y3W/XEjfMCC68jVOLQK0h8lKikFrxUdlkIgg6RUeEW0rXVfDadvhadjJF
OL3ExcBzh+vsj3kQe1jMRLSY5WmrUGjUZ12t+pshU0QrIpA7dH5rzfg87fAfXNoY6TPPuYAexiPr
N85+k4X1mKxyJiau5DveZw0tfJAuPj21hIMAvQNz65fQdEliRIevLRK+9IXz5BCC54QRkpbQRCUa
F9nImaqzCcfKvoKniJJ0VK781Es5bF9fQ1u3NSc7nMZMCKWiG7MAAyt2A+oVXzhWFZmOFEMA4/an
zx5ADqi5eLdXK8wAccFzlraeOxJHydWxYaFRBqFylBE0RPxyWAZFH6vquS3TEEFlUHXEKtA+OKAf
P55f065Pb10si4ycF4XfOsKtKO2eRjlu/rj8S0m1Q4JdCdQel29gLSS/KWNKibmvHcGjRWZHyrsx
kNtcO4MAU4819YUj2aeBb1flBoIezE6zLTFNcrh8CiqruhroFxMuu21BVZtNy2bnDjUItE9RUTbr
OU9yh/DfW5K7Ud6H3eFsSVWqLCuZe1Yq0w9H8JRDmHLHE0v5PMfW1i1gGLh2JyVermgue24Pc27N
3/EGGdTrysC6j1AFZvqzUsGX3Y4UWXDvl/ToKjdVGCvr5ujvYfVqPXwRuBKmmmtn4O5/jmtgvEyV
9tSF42Jf0O1uHU0H9fTV/SL95Pcj+g/YEWOsgOP5TWS6CHvl3ss7WCh+S3mW89O6FzJJuigvaw+A
HrJ1Bd4JyjguURfXJRRvbEhSYLrkEdzUO50rhRHy5Ku2JOHZYY0Vd7NIAeuSA/fMwT1uGRgD2+pP
pBpyKG5KoYbgsfXPxRoOaf0H2Vud6rMi04be8N+5B7oehxMupRRc5lWfuVcThk5zbwm0hF9v0NBi
x+hruqyJob8rcs2ndChyxsDBKCCmHBysyxLvCBoLPC6jwEGnqJKcByddoH8RGnVV0vXfzzauuHNg
gjUYgSJb1hZ6hCOpbbWa8mD3sjILU5jzArnrcQOTcD0oNParUvT8FEir+FpZ4Lbn9KZmiVQK5a0l
9fUxe0SlfPGuECaVuOdq3CxnB3NvKDFuvm0+ir3OmOiUmTJVad/SNFUMJ8WogcewdkyvdnpavBgH
I5NslRqFVnv9fvSjjNh1qbYvzqddS1qAsKPwd5HOU7s6rP/c/ydzDj8y5qBX9ICWSt6TJSBedrn9
Nt8UrjFplmV3U8hJBhN2AHq+i4tuMAXODehu1xrWRYn6fj0G2kNI6mSVCdS9Rw/QumM4B+dTVwG0
U9V6F72fdVj4KJSuC9ve9Lfli+ZKnOaX3DrycMwiSv9YOwxQVBNhYoD0vBzrpaaKwxpb0oNJM76m
HiSc8KLzPZHM2vNrJ+SKmTKAMCBQLO+ng37OuQ/0ltIqh0tOpnAED9PEUgVjgsy28U+loU9a7tQZ
AuCSdWEH7QIfVDE26GmZUx1awVuwTwTSjU648OScDYNdBlawk9+F8+eVz+2/5HxBfcHhO0C+bq+L
LlbdHMFWsKIebp6FXsYAWS5rDFOECYRKOScY/O8/tiOqPvSpBGqjgzS4+2u3E4RsMfcGOD0iUIvT
xb6w+fC69FGGGxfFEcgSj7wJrGFpy8ElI/CCgBzaZlsXDwFxihegTfWeHjCr1tV+2mYk/SWbvYxJ
IzXtZBlGPo+ky6xFX5A1AykYSfY1PtLywpyw2j1QiIodRPQdS48EExKo4x0eS68jkT1gMTXg/Zyq
+Wrbn8UV/1Gz/tgeg5f/6qCIAfotKOHjTiScyfBH6/3dG9mX0irD97f23WWunm9znki5ZjJYfNHY
3NFkeQm4SlSnuI59p9PxY4igk1dJxLud7/In6PEGph8zi0qRQXXEjQLEEY6u2pgx73Bi8xYL3Hs0
BzVOFr1y2HqndC9DAeEv7JF4BBU69J98vifltvC22c17LhxXAdE3IyTXkBIok8lDOLybFHTAdhMX
IwR61CTr5j1Ki+/EWveQt6X1PQUFi080+aaUnsJ636kDSvZJUANnUVKUPb2thr5hXLX7TBMmqzJ6
r0jjTVSYNJt9EfADb6b4qqPR4vCaXRTgDJA+NPUk/Tn3DlmQysUSWfbSD5oI+HAboQQV84xRfiyU
wiug36ZWfblZHbOKa2XP/wf/i/4hT+XW+HVEEUqQ9oYM2DUBj2ZU7TVVfAU8kJwFPUGW3whzlj/O
YCr0t4VZyeBr3qz92FvJOGS77UeMclZUjIRiqiNZD1/ZPESanqn9JQOwtnzGboxBu6wKzgm4V2go
cV1QgjIX/BUxskxB5YWt2EjI02LIMyjLu3llxHhEf1XFbr1kpMef2B3aUxKaRlqvn99EjssHdj6P
f30Uuyo3NN574bF033rsG7Eqo0VQsNK6J/9uHHYSbkQLdGVDV0YvNXDPclKslXykbaMnWRGXfQGv
GTB5juq8RBJLVx4L8JThhdIZrHHibegIsIvQ4rlZWC/r6yo5ThzCM4OWUYs102uWp1/ht/HqOEML
u0N3oRnwof1dj9yjj9eZLVVASv0K6MLJohIrZ0fK6VLydWG0KJKPFphRAJtb7MMRBBEMkQF8MW+W
Gp2DHwSXWQLMf2XdSh06lZOV3vF8+C3FiN814vX68e2E1HiDomJInPYTMUIKTnLjE65tFq1GUnhN
1kk2I7azMPp2G9m2bHHQcXnWojj+CmrXr6zpSPfJNSEDEFXkcjazfXjteTtGJcQxJnMHBVp5Tj/o
HSK1EFl1yoJ+WqvyP6O9MAAOpaWvArDmU2fJIwB86k5MsfDB4OydiefVwy8mzWzamEpQXhoB830A
HkRVCoqVLU7FPVfGPYePYxp69IpE6BUpk0pG5cCNQmtf7NPNwigs2T93FyhfIr8Zp2xJpyYlhn4r
IsKzMxinuYEXKTkC7F3jGg/D+Es4d9K3f4RhKrPLifGaMeWW9GUYv0Pyb3mTse1+ek13jU+dTfVa
Y4ea6i6PI0iVGkw6cxFmQh3QGzSoQVuz8Mh/OOVxTR3czMkGG2U4FdRX113TeZ8LPhqyJyCqeCzi
kEIx86NdJH7uuMjpJ41BcVaU9/sJO4+w83ql+By70yVZMFecJLc+WxiS0Qhmv+I0VOWb6IhnvNkh
z3xR+EsSm8mHhdHM9vMaz8qRE05qI4isucA8vbabDNfD26Y54gKthvpmyq06JMT2xses3Ds7viZw
NTvM5vPdlh+68jCwRq3PEYFfN8NXSO+Nwb5qTqjnekP4pNI721BswGSl12eh8BWPIq3g2TYZI3Vd
xyI22h68Lwit1t8BNh3KYrDBj0z9LhTxF3kLlRTC/FVLw33IYXIbLmy5LGmnyp6uTrmm5HeZdr84
II/r86bnOcDPmL/lZjaQPGi/054i2L8O14o1nxiSCtHHjybNAOpDh3EoP+Qq1njFqj0iiOgYQor8
kLmeKNETXSGp54YQVjVMGdHn3a25YXjRvOA7OnePRJHgqvz257d7UNfZ7D+FmraK6xJsbDHbhDcy
/S5bFxO2C4BQg55zxoBHaeLk6tAFA185t6q2ZQS1vAwAnyXn7Ld8Ox/i02u1lbV+mLX4iw9uWxTd
q/Ct70fl7NHeIdDemw9Lm3jGaa3MMO5NcdVD8Xk2Ko1HDAX5PT+7E/OAewHCCrFwLvmFYLP7tAe9
lE6fnvGWvc2gLNiPrhTm2mjE+FIZX1Ui8RHZAcpY2Kp1XCXbE4qBQXqNEAH9xJD897lQ36lItl+/
hLnmqjHcftCiFKfC6tMy5YTS/aFzyTaIObHk/r4J0lAVJdeXzUMbJn1KTfWdXKaaSiWFFoULCDzW
RhrNKHzXWNtQ1d42akRrq15aUx5lAepy6BIeKftJyXjwnTQBI7tH7NzsvDMTmxi1VPB4yZi8XqPC
tmHZtegcdWCxM205jbKLWztPnzjNtzXmPsUD6nRfu7ubTnwSLHI2tgrklr6EUPQPrrZV5lZVE2ri
Ut7B5stRSQC6Kk31Q9i/DpBiAZ7aLesMZSkWT+X/btpHfVTHqVydwsp5sigAZGKQG+VKabJInsms
61ueMJ0NEjhp1Todr0bMSJcpYI9lsmFIrJ3SvcogO28U4KORzw42QbCW4TFQf5mHy8AKu0je1atu
DAldBJEKCFPKz7XceHEUSOBc8y6PvSpG/I3ZT1VcmzgwtaRce/Tz6vyCs5m+LEeTxMHaXphDFnai
M6GJOJ3CUrZRXOvuJbmxJMguzBHT6l4ytI8EqZfUXgstjXwkhOyHcXxXzecoRzPkdYg2AZjowIaD
02scLSwrxeFaoDz9DMWjgZ5P7pNXruwD8O2URyn3MLVKfmd9V4ySNpHS03yHB/573qJTEdHsoyFh
IzNZCLSmSf4Qs06iuYEVbX2kuBtYVMIniMkCdjmKGP7DZoDg14zgYp20zXFQhWDQm951QkRsSqPB
VQthuWbUfYM6iYX7nItVlgtQHf0SxbTxeieFV3F3ntAMMSZSlsLJ5HcURNB5njAze2sKc8o58bvS
LsZiRpgDxteD3kTOVz7lC4w1YkRlLN97ZJqUxFd1wSykWtMnfY3ip8vTmp7lWRBjkToGaY+g4MhY
LXVWhlLY7+uIZaYE6MFAsqqrttg2EgWkZEA4MbJRcgJ4g3FjRgkjuQqQwxaRXjdUXdZFWdKZLZVz
hf/Na4/cqShxXiZV471gmueswEaxqf8/k3r7Y1WG1YitmW17fVaj+7Wm0udEgH9sDxGhkrdk0yGq
N6XhY3LB7msRsP2/z7W1eI8O2nnrL5Iw6wox1HXv+AZqbIcBXVN4SQehJs2M4BxCSuhsdxENorUf
0Ai6CQTfC6a3aOABOtdfkfcQMGa9+GbJ6E2uLAfwkbbVmiKmg+71kUifdO8LEC478bfe42dwqwT6
GK0kXnNPn18xMCSz3TN4oQ4SvySKqzo/ubT6xEGQ0fxc6bCBa2854fDeT/xoxKdVX/PaPZiD2vIF
S4skbrFnTAv8cysYQ2r0cOQ47FwvxJcBWNv0rwyMMKn6JCKfnhevV7ztrJ6Cl2h/acZgA86m746Z
FMU5d2OkgE7xuKnt99BN4m/hce+hyGsJWhlAatI25fTu2EDYvZrwZOpgecBsUfImno0D5ndmx3rs
Q586R8EcwcoH2mQMPgmIZhN9If7O1d0H4k/YPZ+7mAaJDPARp9xFsFyhJRf4g7ue0JNc72S5tvoT
KlSYsyZdea+qkY6B9pqfzIe2eIGjYDuDnyeYl0sD6M0TqEJBSq2ldwEJAynul32fcW8kiMG9cWO+
mIfQJToaw3vgWwEvS/UuCbzMN1zQshLH+5w+lZfx9PPLFys/rTQSfUPuYy35KkW+OkQh9EcycbPW
FpxwuAh44r9XQ6k8/tE9447meL2AYQoKFByEXu3MouuPhw/uuZx/QMEFzZHYzMfqjkGsXUmLdnI3
6tQg7pQ0lMQv0mWj8BgjgXrRtvxXr/O1CFtn0KZHgVUZdM+g/FYBrfwREB8GGKzusffHaiEC2Egy
t+FP7E5bnSOIfTsxEU4hl6sVcfZ0VzjFKwvgZ1SsYB+oEBXR+k2DVyv7HV8doBXwsEfNshGBdmZg
offvzv1zgaIib64dOV9LKeLEAyWwXavEp+2Vp8SRkREWQQ1FdpEne7mgbxFZUd7pfNdkdxCtc8OI
DV/vrziksoOcXxpKTTbKA5v23qLtIwHb6KEEFM2nc+/VV1FWp+0I9kG3vN/FHqvWxffqs7gwZzf1
SKKCd5Em4OjGI2HLJZ4ZKKUIwlDc+rwI65fNdPMUsTjXTUD19M6g7aTXFHWeftYBEZHkSsjE86bo
Lu8935Dc/5hta97tAFW69gBwF5m9BHMYhP+7zGQYHJTvbOwXD7Ea6F/nvNw4HriT/+bOIqdqioyU
qcvEAPZl1DPtnbWkK7Ok/UMNukJk85mFf4Xw2B+nAVf47mfax19AyoJdYcWQzHFJcV3R4k2dH3Bj
xc0GrX/tI3lckHxbJjW83JWi1GJUjgh32STzVRIxbD9soYyCLmVaBga35a9hXtKRx1ovD0Xmskj+
lLbDRg8eCkd6ud5/pV29E6ocePESm82jW/FKwHIzoAtRioJH/j2IETKQwAmCGsZClN+u64yy9HQB
dyvaqnyy2F+BuldX72SVPm5ytV6GOro55u/uDWYkGAyZAg0gPlz32GNz/HmPK8sbNV2bv2s2IEfg
Nk+952BJAwDGACupUADUg/dqlvOhmSsq13Zpbme1SfavQ3jGpV1LbjuuuLRKNLfsRChGLIXTtswM
vF2Otgpk01HoOVm/gdxu9lxJDwqyTj/t88t6p/+wjXLFg+oEWL6ugF2kVC6JNa532/nuyftvqYeW
hSBAoaCA0wkjBaCvduYbpU/ZeW9I1feRD4JpeNQAbDQYZDbJ3SRm2Vr7JUzp4o3scqSKqdgd/oV8
o5s0SsxoSNFBseMF/D99VwK9qshZ2fqrmaYqX4MKjxC+G8Epj4xAHYSCoyXuzrag1Os4yLTt0js6
GX8ac57Us9+3JgGQCshDCsrDh06wZxTUCvc784qq8jy6l/7IA72FAWU/mV0FidEakE85OJia7NgW
k1SI816WuOMQHW+T9zdw8D94gPNX3s292tCVKYOLKPLcC5472NbWeLm390ApuNhNOmq49kqQI2Lg
UtKewneqYmDz8LU7uf/6kWHTBySzJa+yRQ4xuKeWa/W7huTnf1WP/J/pGWz1ZslMLZ61K7p7eiiI
Myb4fKRaVKfopwm7lU3VNUm6fmFybAV9DPcSHVX+vTMP4CrGhnX5gpTDYaYSQkhajcfGTyzOj5Lu
ui2lN3mj+weT3nNlSJ9gm9wYyQVhCww3Y/G+l79vfk6c/poABfgEFP2YJObEV/ul/GqRMhF6L1+F
oBG5QJIYlPDnt6L0JxudxTLBYWB5mx/8OzN4qfjHZuflZZn15Qtx7LdkwP1w0U0WbJspqPGkXh6U
v5voK8nKVZXltF7SO/qgCiT3j5u8yk1YVdDoLpZcQhrROzvukcx6skhniYEZMTdaIac/zUKBZVL1
GsIjYvWkMi8oeU+kTxOdkeFSZzyyq1hmf1SzYBiGLlLbUPHtkfkR7rbAxrgWEI1JT+T/kjac/fdh
ywOOLsqnJ4VuJgT4cKCYfFAOKTvF/gPwy6CA1Cpa7IxOmqQCvGg+sRQ1AVWmGl+VqxGkkDUBc3PY
Kob12KAzP2qVFYOkowsAYHscfUilUTfVQQHWmB7tYala09kOSoQMYqVTRI/fNAydgFIdnwBUCXdK
aglqFG4ApLe8RTXwhCPE0qhl4m2zFnOtH3UTYujKYdwLWxATNRfcRm+irfpLo2J83rOHpWu4WSeR
o02jDFjgQFkuLZfC4i5B4K/XZmwoX7L3IDLwNtP+TOuI/WlClVEb0jf4zhWPMd/vGa1d87bzYVqJ
5SFNWJJnLTr5YfsvJgeEbzSsuiUWOvrFPtjM7Ts772D/7prZnOWXEgM2pFgvZJmeJ0k+Pd5MB8Gs
mHmhNyfd12euiT0rScCFRa4wNvrMbXrtH6I1VWi3dKd4tQ4Oi88JOtQS0rVd2lYavH4gZyRjpRkg
qLctCNr5jxrPqozSLwk8fFcrCXrHUgOxvmyshhNbRmAcWAJ/qqJTZQGQVkGPXiHCSxc2FyFO6MFe
zKVx8KrWarf06FLzhSGkSVLTrPOlBbz2oGPRzYVQc+m0HvjbnieqE/sThxPlABwjU2d5nF9p5Dng
53nf9pUbOfLYiaIhwau8oo7IPspT3iTEHx4ZHkxFdSZWh8wERjoQLUuvF/zEqlPh81MqAkVFrOQP
K42IUYZjN9sAbPu/SdCi6B0Wy70QiRQFatKQKyd57sjSR5bNX8nVsgtTmPc7kVt2S5M9dBANXGfS
g5s/3gquDvDl1ICwIt9d03RFy/SNextBt8vbnRpCq4wySWf9TEBigY6ct/eaVALxKVj/y7E4yNYC
Ybg4wcHRo/cqDlkZQIAzwiDhlIWyfYj4sFckVb6bgm8oWgur9aD/442OEym4oDeIkz4jOTKxf1cu
qfe/cS0PSv0KqZOeskxfYbNbiWJCcsQBpiSD4hJAQxQ+tqOQ+bhUBBqDMgaxJTixU84Xsn5qmGEa
Fx+AUmyM84mXWp1ursQdAsD3kTZS0loFy6hVufMOvBVe57EKdTq1v2dwDG8BvAIOk84ye6MsDUYb
Tm4kw/8Rh4CRMY6LEPDcGl5pAFEl9VKRP7zv7J1OP4lRgE58I+lnwSohJ/FdeJ1/nPSptp/wSzI1
8DvB1vsCQsgJSSBRnc4tpjcRUaVkRtuY7+mMBCO6F5AlPtGYvNoRTXkzJFEJjwYnoTJ1yvFj1TxO
FS1b/6BMStLR4rkfCcGcK1Geg2V/rvmehZhM7PALct5TsRXp8kdaoXFgHgUygO4Ggno2VjmC5+7c
zGuR3xSm5vgmIrSji66n/XQEuve+ZIeuvLmsm4v9r7yvjCxPYIkyMsULB1fV5uwxV+nPbw/8LCPp
NaqKxcrKFf1Z2YnfZKQfe0pXyasOI9QiVpFH3IkPJEN/GSF96n3Iet049Juf90LuLK1E6S15blRR
bJrAhr59gB+DRhjVUErvOR3oQ73hAU3AaKsfmr1Bvy54yOm1aUTqjXQ1tdgZJ2YtHqbhtWflLjUo
bRiXQoIZvOcTduf2Ij/NhPsIjo7OBZJww2TjglrmqufZJGkDxNVRwuM2PSX78MXfXkAP8/o2RzxA
ddrH4HOVJCaXCLcm5N0tlL7CBtDFLtsDguCKYTW6KNjW1sxo72mQbkM0/wVDxhm5Kx2ynlLa6wzm
7UFQ8KiYhL0M8BHWOzDn6qvegV1fyyHy0fVICi4c2Av1VYTLc51POlT9n1B9q04RaDsvmKjD/MlA
L4y70Vf9+1tX9BqP7dpvk/Em+HUGY7FMicUuY3s3uaQiq/7SgI6+PBADRWMpWxvRAUuBJcLd7+IV
FhdZXAexrs4paBEjZuhPpERVcmPwmN5MmKTBbCm3Isc/6P2IsLnxrUnodqBGomaAUYKL3wcx3/7x
jcR0POQ82FiWVAnBT/ljENCYM7tmaK3K7AnlpnAIlFG713Ptl1OYkQf53z2TREolV4UYhP32ptCU
xnORJoMK9qu6Xh1AMv5rJ9RSRBWYygNTflrZiG1zaZ/IWGuG2NdAwQaQO23wgQoAf1tyy3h7F4RB
uHK50ZKDSVrbPnXvo6xIeULh7H7/AqtX9duRRm1kuR3IInq7/iulZOXEJmCwRdzXzpDLcUqLmKA9
Ucde2jWIZsH+1/ru91GbcAyhFP30/2dLaVtrO2pstNtbrV7iTK7BKtCr1mbXssTCJYy2SseJBYNB
TbX3EFGJ8wUSucVH8PuKGdgC5cSHLqlnzSMxBQKKdMKi73JRHNPyx4hcOPi/oj4apV5+eCCW84wr
8OmqWKYQXrnBRFM81dhI//Y8CdH3eG1o5BeUSaS1OBXzoMXy+jmkeJgwivkiuU8gSfujeiYYdvTf
HCo9RTNp8bik/98u+xN4wDEYbrsce5nGlBrEFtNi9AQWFmv4wtvCjQGskb9mJ+ka3cHssxKxA5JF
eyQYCWBmxQ0V9yYqFStmC0R+hlxA/gglZIFmZ2FzWKPV2U5DfJayHMya+quQBxl+m89mQFTq4Kll
mQjpipZ9AluNBXFOaxxqi4qY0df2hsN11gAjlOi5r2bdnJgkGORe2CQrI+ZzuO8HkwSmwnRsynai
xuyynQm287IBanH8BVttpe0dpPG+SeQ/RD1Our+6wobCsSvON+TzV6Nm3uwkhY9g7a5YWsPGhRaH
YAcoKN0T1v+WgHw/p8K4j/O8GLJ0rLStl4FZiFbYRw6kz5XH0frxRK+nuP0rnIGADemd8t2UWYxN
bAdB/wdeEsu5YwoWqpfAGroH7f3s1+LB0xXedMPjNcww5fCGUoJ5JQmsJzvvKIvK+EXSENhyt7EU
Ww72rPWTmAt7iZmWC3gIeUvjNu7k9GaQEIsZSj6SyRqj6wAwQpoMYBD0ywfrlVnUeb7xvWa9SNRB
ZHbjpzN0U8Cnqlr3DSLSvB7bb2vvoCJWzU2SQhbYB1r0YJnE+KMT5uQ6K+NfKa7ZBVA9nROPNYWi
o4NPyHXC8aNOsvyRFaqt6F+B5SGzuGA0iUbKmjBwOnfOByeAEMPTffA/gqB4BI69UD5UPjFPqJYg
NaAalG9HCoeEeMHPTkZlrZNOamyh8sdBqMIfiScXw0W3Tu3kUgLoZsjdgC+a7ym3KEiGEydfulNR
RmXHHW91YCygx6oS5R6wsyx+OtBZzpKgZ416BCJKkKS6N7/o9gwrQAqB5khDrycbnA+b1dZD9aQo
vf8MAd8ARYabgvw/KFBodgMNAxn6xUWDZbQ6gfGZhmd3q3geHk7I8Q5ve6WPMpUwAWppyHsm9nzy
wbM/ETQTOKbg7K+gm01jF1bNyukCWt8nIo7Ss10sajcv1GgUZQgo1eJ13H2VoT4QxISZfFUoAJlG
2v78kAhk1d3nhxr96ILBHR9lTDMTNLmzCTO/ce/fLajeM3S3QEfScpSHnseXkBy+e06w+s9ezVwm
yMxfjZAQuCidBZKsTprAYRLZzpWoRZ8Oi5UciV7pziyA7QOjAXdgovte4CVlflaqwfyFe2lL2nOL
vxl3oot5rUR5z69thcteR5FUaTOG2f4X8j1tEAhIC+7ZSvsTDxklkDZ2zvTU99OKxGNUzXDUrcKq
gd3UBGQj9HYcjmHtrMa5XMtSxPalOrzQR7dEq8QFWThoYEeWsKTIoL0OlHGYXdnB39HufhKuLp+S
oEA6MrH3/vDowIGl3CXUGfL2mUR93HrKOfk0yTFS85ZcdBhyk7yPYhsn+C9SkKjFqWeKa1ibQQ0H
a7oovssyXrp0La9/UDbWLrqRMixL3PFqjfqW/JsPFuxciHxidNPVaVZ0dU6jnT8VjdxrPirlMfLF
eYKOEUAILGLEQ7vTQgPRowMegzTO9CeVPodepNl34T8ItLNoVxcNiP/cVxjiAoNfc0XrEXQugxQM
02gG2UtuOE0qqe/dedMwHr85p29ly6fqDesq7fccOPiK6mmHbsE81mxcj/h27XgALvg9dRxWna22
oUr58XDicVibAHrMIXaqGW+jerSzbAKzFQ6aFd3uYV/5nxmLdpBhU6eqzWVz1WuzEvYXHHjJgRCT
cFmw0EW3vp4O3QM2XrzZ7gWYUBlXuB2gDVOo25N3RoiAlfa7/+rzPwRbWx4Z/G8z3/eTedGyXjGu
sXVsnGo+yTwGTs/r0Z/NZzWQheh5IWJcR3jkE9BnahelDlc1Gr91oahJzF5hwXTHGjKY96XLaIDe
X0KaNxTwDz78qvJO4N5txIkwinngFCyxF/hTiBd18BrlxDMQQQIOhPQIeYOa2m3+nto62c+7J33U
xRnRThgBDvogdhwm5VYM42sULt9CBtZuFowep8jRUl0ztYhKjWXTEJ2eblA95yEj2ceAjPRv+6Ee
/NLXxxUKnAm4pWhSZEsqDdrL8Mjbv+cmVkiYAD7KO8E3FZIogEl5TdE4T/UMGAUJjEsfvuVtb9sB
Oha/Y5yERAUeI49s69juioBhKvRlaboIUbHPmuOsR1AI6p6WE/Llfkdhb+aQAQle7KeHCSV/nRh6
FdM26Z1YLAMQcWLAIQVulGSludZOY+ubvMryHCnx117YOLMyaWGy38uJtXDYZD/hSBhNorH7IuaA
3qZWSmM2jH51DkH3FsoieinfOoBIS/F0FUBRHSX/w65Wkk6cYL/S+ZmkPlYuV5PSuPztbXs5fjSZ
V/Sou6kq5qmEjYR7aVFlHPsJ20ETc5uGHUH1gGZ79uvAtsJZyZ/2XcBcbZ8F544JjqLDcWGXQs3g
ZL6jF/EUPb3knXxH5AMe6qgXsRJJUOCus4DRWmAObPrg8ZX1ts/MbbnyGnjGxmWWYOTFS3zKP4oI
yFOJvM/NzA9VJqNvgHMSi439qVHxTFlQP8Fj/ekSNKKk2/6CSFrEIgytxHvqtMI0pdbi2ny5vhFR
qaUTno+jwZ7S5ZCwFX4ArUs5uYuij2MDfRYPM1le77TWMdSETHbCttw9JhzEFM04OS4ayS2gdzcf
QwSfEIJU/XmNBZ7UttW5ROxTVh4HB/JVUGTqAK3vSfuoQ0r+EOOJxOGi/RJr+7xuaIifPPi4t4NG
hduIW//xRcHMr/HZbdNce2YmwVa7w1B6tqUycSE1xJvo/ciCMxvB/3wFiK/bUcsBZKhuRQgj8UPf
IA7gyEzH/uy/LV5Gk1G6AsQVr4TTaGNsnviaJ1YE4zCjlCiDDmYXU9r0CHj9iNfr18GoC6/7TeYd
HI+WhtsDgw6Cz/ehHj6Nx1HNKySBi8mtQD4pMvNpGsuvghbV6WWi7CV26NCE/ezDOwNfDbiTHmDs
LPQ/y0Y8fju/phTyWyJ/tzESxfkjI70IcYm3fCJmBVWOUpKFNXSEcUvp2IHCIUqM4/6DO+P8EyU7
E7KhSGAXT5XxcnNly1mH/UeIrHAbpNSUZia9kxh0GlkGsIuQ1nqGjzMFfsOvI2ecZ+SeK7C5CFCj
JiYr0OhJ8A+XA7fqRd/MQDd/hvvrvJ1p24JWBwPmJ6nnuEWoSQcDtfxsgFLiNjrO22ecWYsobLuk
AxiH5aKr/qR7NoB4EYto3m8VCkun8T8JXGcuskesOxorX1+TWHAaSwCogOkYZzqFR9SSRAlKc5rA
Qu9YkiKmLuKLCn9/1yJYm1E7h7WKeHsVu0o2Gl+F0M+HBc3/xCR8Xo3JsZZQj2GOzIHPMjMMAmNI
vg6IsIs0SpYF4yLM7Z8OHUaQi4LxxLNr/zZELn4jYH40pKw59IfHfrkYC4gKlQef8ebx0SodZ2mP
XntUSLxJjR8l+PSKevVlgH8+NFvcJ3z9F3GUffAhiuJKk2F/WlKmpZISwcn7HHGYCIYoQplTlsuk
Am+9s0fObT2VN0h0DDU8OptGUv8OEfWlrWryQg5thnD7wF92tKYUEaRafZkW2dWLGeseSVVS8U4S
dBmdQWoFtNbOIA5Od/p4bDZYxKw3pqjs8/8GnriSHCOJuxSY+5cHR1+zj8GWSSAar3E+0daKONfw
XnioLPkT/QXS/8UQ8BGKOYQA1rSHRmiJQH/5ZKpwqHdJ4kGyg2RwiafLh2XUw+XaQgJK9H56wKXo
1SmWY3zv80V4OCU5eFi4RCWTd20IrKhoJk+a0DWKupuHucKhA1I3MlBBMvFFzW/3IKqtlfMNYjUL
HXilA7HGCu2Fb+2PIzjwhrTFAdyDHSRNuElPblDTiNxKMKOBQ7ulmqbBv0xwCQEsvVt283eqBpVD
ZQENIyEADuqjjVdmY6ponBR4x/SbzI4VZsRdlhMXIZtjnGVtN3EkizX5+MOBL4A7WpUQrPFzty2J
RqrGUsfDeeLyxvX9D5OKc4D5adX1enZJSY0e21AU6129WdB/otJJVCIBRRkRBr3/rpaN1MVQzyqS
N+NXxKCXoaoiPIxnueAmCmiunw9/jJPiLoQXoEwmHXxa++QCjTVsnPETx9ZAxisCFDfAZE9qLOV0
3vy0a1991o/MgKXzd2+2eQ8k8+UaruxoOQ092hi+f+O2vPj6nJ+nCm9avTN3JggCWnVl4Nh3U77C
UfUvgUauQ0/Q6FAsbDPmMCZreB5hy4Rhme9/4cXtjUT4CpQQ+XH3Z8OqAEUxiU6703MgSeFBMSKK
h04OASeqQHJ9th/RM3M+jT1ht4YAJteog2qCd+cFMHDq+qp6N6x8q4D0V0oV2a3IYMDlFw+7Lpux
ZIYuQauEPQv5VnLUJcHtlgTMX318oXl/b7AHaRGdnzvprkIK7hVdRXrquLUiiGC3yzM23bIlx+2D
5sAONDkRX13EXE5+0PzxGBgwWrszd4f0pFmWxnpHmuveFF1Ss0JXWzCFyv198RLae78ErkXdR7qh
bZ/t+7oCHH7A+IQO5JNWVcQ3MiSXeDti3NxLy84Dqh0yX2BdIgLhImx6AZP5i4DZJ8Q//Uxx4Z8r
kWSzu4mk0J1WVfsRST635LIyrBM5yUkB/uIbxtDWSqie7RVNgEvAVFDm+bFlIz3PNTVwbkNQz2qO
E1u5K37mGWUDlgKaSpVvFwYexSrWK18NIS2eO2bKesvmlK1GjoSTzAgB/+MojXlSThGz0QB23yXE
xd9bl3b5H/X8/s07Z7DTOYW62pH1BBuvSonsuSyq+lU+L1Ct7CJnM9UK2vyEuQHZwz8XAQkSXKjc
hYXTghHc0Toe1KhiAQVfUE8wx7o8DO6SLuhWL6LoX37pfnbJVcw6JTdzfPtdoIE61HOMJDgXWl6r
kaUrrFoFTtGFl56aRaSXx7C+mLRyt66UyU/6kVik9czIlxOhR1SMG6dsPU5hxXrzih8BwWOO1uyc
5DhNWH4ahxppRUpcMEHBPMq/47D2qXCU2oDUKeL2J5RruU3lUDFpKTPdZVJSUg+PqQIw705pGgEB
lnfV+YAT9Pw2PRvUicMHGvN12I1B1x4+ZOwTk5UbAbZjtG9JBU4r4e+KVbG0vdliBVh1JAGhnGbw
TrMasLuQCuquWqGX92fYRgRvPBnZEC2IHrqt2dk2ryo7GWrVwrICh6eKU/zPJGixbvMwtSLMsXCS
kR3jp1KFocACGsywj+1VyiTvvCIhfOyKWt6GKYUM3hh3Y9YC1EI1HDQC13PWY06OS6tG63e8UwBG
rhlsHPYafDYxuuAKUKfmrDqyWUnncbYt6BHL2q2jS6noilYRUQJ80GHr2Yg2PWhCfD8p3aaPW00o
L/9qP22a8Fy+MEOS68XHAVnHnwN53Grdg7zymQ1/bTk40rldquLlbtGiHl2frQsmAl+0PSjUUePh
mBTxQIQjGnB3ShX16bPEdEiy76tR5SMiQ2GoUlcsCdis6/U2kRBt+FU+f9qhuZD9bhY1kDyM2H9C
X/cJxcrZL1z48w7uxOz5hxqyu3DCYpfRadozfph98iJJFXThjYIyfWC48TITNxo2d+TEFFYGa/5t
QqbhAzFGqhEKDXaxhZve4qa6r3qNpwqEG1DK/v4Ymf3MzeNj5yP4JQEtO5ZQAkG8rJ8ASiPwssST
oPgvCFziFRNQd1xLuslGECt5D09REjlzbIe1Eo5bgtLwF9tQLCmN0sjBQk2MQIEoFvABpPk1xvDX
mRYn/0iVqXkN2bn0sffvwocUYxg88fwS0YERsLpx2ZNSj6kc9g8bKf+Wzw8XiIkbih4XTpekRnsN
lr5bBn1zwmabdPKwd8SvxYSWMWukxvnQkYN8I+AFkIldT8pbCsLr1SE2Baa21yU7yEsas5NmFW7+
OrwWj5YXIM/kB2+2nICGwWtvaSn/lp6hIyBCaJTqH1fMvByQWKfngXM3kQRkzLZmSsi0aF6EyeJe
JHBmsokGPwage12+SmqzxC6e7y/7EQXrte0uyCw2LjSQkQrETZcOLFyCbca/NWt9IKLHVdUISjyb
5pF/MykhUmx/dR6HuiLjaC8PFffNYNudcCv/W0TsHrATCu9lH6zD9JLPW53/V+fIO/z0/trX90YM
L+N75/YVqwTBCkiuNoMOg3t5AsicEK5LFc9rITrpiewaEP5Lrbsu9KH8rDY2TTW1Ec1TiCtW3Kfx
6Yp8blilC8E733r1N/ckPqxmj0MFV1DsnRoc02FbTau7/4WaxxEIdCzRpWJ5w/d6XqKHze2SrRN8
3ivvxH/pH1OanbkkTCD/NE2UMSXzSQxNWltDLO8ikZyW/w+h1GWMVppicf1px+w7q43NMOBAcqEM
YbA9ZpxAjNwkFvcgpytcm8+jxNSzMrHEJvP+AfWdgt5uJ6pKiQ22Xxdkb1FGMaqVan54drmbu4lp
3S1+gAmkgFD+Jp1vH5UQInTvFPcBQG9kVZRUfqDGOYXd4S81eYPzVd6x4yULL8q4LhBMgqgY8/bz
SkvkaaNi1vU+v5CWk3Y8UE6frwbhsCGjY7ZziTt9rnTveqokpoIfCyvuUJbRMDAnEjDkcKmjqVZu
AZHQgSW1f85AcwQ165Hp+2M0VPOh0L9ZjhBgHV9cuA2ckOhKdmZrfrONeAnbs0fuu7kx61bJR3mn
XB+dGgdpTeyeDmeeEUAlPTMI+taUFMBFXieqW3cCwl0uoH71BbtTDGWKzsddXVakVtznnKZnMogV
b38++r0ZPuzwkrbanLwTrIoMcJ2I3HfWggagDMaDDfgzOnC4KkTOdNFiw02xsdGCQnG3by6HVjqf
hkjxW8TYl9VlxMDPHXsNfVcs3ry1RlrUwXsSPz9knCHS+RZqEHwjG0SXLOHaDtYq8lG1b3zUbpuU
/fO5ENdigpKwEy1SMA/VHOG0d55aafhSo2pSoKp6QRugyZwdhvtkHyMrNdsURPsATbVfqtEehcO0
qxd4f5KQ9QbvhEEOFUmiP9AAcL8+LkGw6y45OU4afJq+yl6FtZGbaFpK6IX6jvpzlLacrNwrvfit
ADado2sYi32QwL7D32yL8u37QACai+nN95IgHPhfo1p8yXEg+zrVeolV07Zms4lipJVvYKK87U9v
0yrgXmQDXt2PHHzNt42twlleWadJjCgSLdjmD72yFfewufkUY7QI2/xQ+k0/VT1kEDQvktxDVwj5
ciK6DQB5YHXHjjHNNKr7ST5IIeQYLj140l0dOPOPRIEP8iD7i3Sb5sN7S8U9tD8A4Pfm99auq1Z4
qJSCEO6jFhycb/rfZqKzBYeHfyn4nk+lSQOqqNmM3JGVb7uKZ/GNveQQnf+5zMDfJLbd2/PQsEgC
z/y3GWiUR7nO06OXfpbQQ3yXKI2w/SzSoNCteozUDcdlNp34IXAoo3jx9v9k9pzXOBfxUiX9i0FH
Wgfrovfk1k8b4Zg+PPs5XHPkqlRQHlSIF9Xu93DF1a3TQcolpSuAopp+YZzwOUYbnV9r5KgSjWvy
fog2dsFdb+eMcSI94J11JEiemZQXX+lArdQUR0WGJzcKbrBQ0Fj+DiYitOew8rZCbWMUPw8VaurA
SON5y0CJ5IgIM8rNuHFdsD7VIN4zZOfF0TpXNwsGsp3dE0B0oq34SkxG5LRjk9iciWnrjb5t+3Hs
z8pM9R/qB0Wb+T2m/2ZwGYnm5pGN7dF6xvyQa6od62mZtnJzYnVnDst/DeoyO3/IXhUvv79QWdwU
vaJu9G+9RB84BQGCqMbt6rrwpt5/goW4gsmixkmiJvcqIR3NvLgGCRaxg5UOSReYNlfpIifJBoOC
lf6R5LCZ4h6TYtTaUijyU2c1/Gmpivz7kCphey/oTO/VAp9Wsg4Sho6BXjIe9jnxfPZLqAl9+amS
9YI8GTtPruGFMQKkzinMcl4LNCuJqHPod8injKrU1UgO50tx7+EmBWhWv7wt3Inp9+BdoQLipdF+
eIW5a/zi8Y7PZH2XTNbTo941nVpoJywI3e5GlhHiimHhX7YP9amHsiwGBzITPekyNm+8+XfiLJN3
HiPx0Em9gA6CR7i9o8rpKdMHubLhcUsEg5SoxDFf4JFRE+3PD2eP/THrUUUHTbg82tk9r5cJCZp5
jkMakmncWv9fo0IntRr0Nj/qUNnzAg76jmJLRJwV0SznIbVluHPHF+OUX5lj/VQMrfC0rP+pgz5J
hv9HKx742IGrFp8FxwNrNMD66KscoHsdnwcsgZ7Y7FSpi9jjT4KEfE17V5VB7uKfOvM/dDzNVfRS
N7Q7lV64xR/LIyEyNsLNYrUtBM3DCYAst8NZV5fMgunaJqaSDZ0lQsjlJNwJVSheRN/9Q2odUms1
NzK47RyDGW94RJd3nVAOVxEiHY4577+OhFEJaa60mEfC6ays+J6oUZIHpOWHYMaXwHL40U8b5Irk
FdESDhtVp9dkhiUeDw29xQtbdtIXdHYakelQZ9M2jdoT2QSJndYwO67wYCTxuSsfW88cBG4BScTY
i88ueGN3BmdO26kwm9JMHxWJiohbvwoXNpoxDTzXhLhGa4qZRWD2n1cWu18qQVsfBmlZYzJubbuo
7vypnsslyVbaCRy0c1v0E+iqaYv/aT7pze0vI4Y32Mq3jjpi8RC4dbgqGpIRSnjQd1c2+c6/yMrr
iE+Hzzienjvs7NhSwnrJIU6XDJCxQhKYJleA6WHYrIClEmJPWVKN3ExpcOXxAHQrbb6XR1Uiqnwj
eh+cI2NpqoNl/rnjzGhBATqIUmyb/pLYOC3CAzQYReaJz2AMYXCGPeLPCoRtpFgBgukUybap3ZV5
iOAoVlRZhPX/6sRAbd8nMau5NzZo8ohibsDVVdn9JVtuB1o07lTeAHxyn3SQSa2w0nid1fsIIqqZ
Rtr5UAxDNBeAyO3o47pOqxK5macvKB6UEAQQPoD3+iKvd9D4cZNoxkuGnsCMMrdieV8zN205FNpe
Bj4SHaHEcsaPlkcGqtaB1VXTTeR3I3BPb7objq5FGiSdYxxPJDVEEW4yTMKovFBjivHHNO7vll1t
YK2MIy33+mUcihuvkgVaNKJIaIEw3dyiJCvto2Zg6J1Zy/ECc2pn1scwJHzVgEyT6RKL1lLiKByA
F6vPBLN/dgUv2SvKOnnxRESSE/1BvdrIpCQUuHu2dCvqTGW0guhgnENyurrmAfYQEAuOBAHcLJ5U
mbZNJSAHwqqvb8n6D/gPOsSZNe4pNSfrN3czT5PXdMgOSNe1nuUEs1shYHmtnXa8cQmGkSiyy60K
rVjEPhtV2HsoolM5CcE+zSQyPLYcIbdtWpaO16947eDAlNEiqKmWvLlZTPKZadTy7Uod6OO4OYfY
zXF9lm5yvwrYd+OGYvozx5RneCzjL5B/tKonwZ9EDjYpIrlaYACUen1bGUl1JAxQ7Q5hsD0HCkz8
mgbqey30CerjqQv/mWM1lEGngKAGsv7G5GU1LWJ0BPFLFWXYhUr5E9ixilE+iNWGuZ8hzni+oEiP
uGj7ZQOFxpGePGLmzhtg09NpsLfkD65SdQ4/wOq6rKWhJOcuglC2+cX+5kspU9yGtVZl5+8m1dpn
e1wkGJ3tieoC58jOVzcYg3mA1aS5m5hqzlxx4K7IT+I6kBTYoRdyv1rbc0nAADRySJmJhtu8V5bo
FV3bNA4EXbZ6chObuMTsZVrSKabl39/IDpXqsvwppcrRsUON2CGeobMtASgq8zJvr86OXpjc5qQs
yzx0MwOSjW0kcUPbG68ZlJhkByDHNJvIwWuU7SxKMg75k8fVfbrWSigBU51oGQIJVmEL9+QeskV4
7mEBnlaAW4J73oj/iDO6nl7UgqDibzem3GmGtG4yQpOwFpyKDjw5O4OoDAVX30mwGIreCXOHFeaf
mR748HPdpzk5Mnl5KZyNfgHMGpzdyeE+ntc1uTojoQT7Iq/I9mlY56lMe4B+FfknKgR8fj107i3o
2fxmV7oOpenSkmxtJgiNrx3iTDF4wvE0AGKwo+i9esqn+UM6gjodGTRX4f19rbQUoP01NMfHgdCS
tZEnr164+EC10rleTI1WNrCJkRjUfSWOPMmr3r9+YTBC3hxnPakVt0Wd+ySXKO+VB0tvN3o0MNVU
zYdwXpA+zoXjWeLBmWw+wipYNp+v5k9C5cERtPryh2dh0j7SI0W4SX1zpmfm/gVuxlXfqbh0tDjk
uFOSANxwOhx9YUYsJN0aGbQvt++czNTff+qjNRWzLI/07D9bmSsH+5Jf4dJwecl3dYiOmKBRO8HD
sZOLiS60OWdmSdqNHom7VI8KwPGup9Kgyp975VzScZjOaDPknZt8NVv9ngDis4oxpFp7LZnen4Ve
shwTnV17fmykDu6jrKdp63jUwYPCT2SjHnaVaJd1I45lhRpKmkaqap8FOZ6VuZeZjyjJu3Tu/xP4
1wmjJAh18cugV1V3phFahImgcoWZaZIi4pAageIUzSDVVobH9AeuQbgzHtI3moZVQS+uV2Fsvr0D
v6QkA3mljyfsOqTbDmf/dBowLrcOuAXLTaOuk7Yj5s/R5KK8CCrzWQGLAkjMSIyoL2NNzjfk/MUP
jXmIG+QrZUiQXM1x0jmoRsXQbWZwA4V6Aee9MgqoGIXJgJ6pu6KJ4Rv1dnCdWa5MyxACoRQHGYdk
1Cfz0T3Heqz7ZagIoPeyLtafH3SoyAVFN3jtmdsk8Q4YhvnB6EnY2mpbt6m7hkWthykO2pU5w4KG
Yd1O19xF8wk2w7Y71g8MKc5mbAQsSlB4OkxTHbeN3kBXsyghKScy21GWhiX8JSxhULZZQfTABYsd
LYY3dvY4kBgD+7JWyy1NAKPAlLF8fuhnOo0AQlk0KCwukJ09A35gdcwycArzGmjQiQLsZ3ncPbaC
E4So+YEcIIaxcPustuWd3z8J3+W+HWFToqYg4XEspYXs3SrYUFpBa6ST1n8+dAIkcAkmQbZg0L3C
PuBSVjOAgq0z4nxBUN16jvpDqVYMCKkV/4cYcdhdg76s0aHbZWTOp3ewVJQK/t6Y8KKfo7kOEZgQ
OHnv6lsQkyYp1W3PYesfB3HhysshZ2e8bbA5zCWMvejAj+NHiJ+MGhfiOKlAmPiLOk0al4Vi6Os0
DcyWOfOmR2H9MVbwYxnqhOve/TqKiohQ2meto8m9Fqov3lceB1l0tzTImM3c6FpFV4LN18WeOgEP
NGIGM6kgeuejMLCBizsZf4PGUbH2lYoSoQvLsHcQr9xuUcaJ0OULaZwN+cGXUqxXSqNEwmTNjb/1
eBjIkslTJg5bmaqhVgX6U9ipaWpa4+2MC1/v4yH9xU+5xnhytgCWFCzkqtvKCmqZoiqRc62Y0R3j
GcoY9UQGiqCTF7XzRJ3N83IwJmzPZpyDDkMoMVa34Y2Cda+e7zuO3sntt9YoUu4LkESoz8frbJa7
fKjSHbRvRuLNsaPP7dFchpyI9i3R1SQIs4krnF+h33dBKX0vUvrBiWc+nwo1xd4GvENsd8jDbChi
Ni493ccAUmOKSIcHLDQQiGseUxHQ+DWfKNn7Gt2DDTD3BgqIWOTiFEuygAyy32u+97h/D2SnPMPK
ITZUyxpYBjOaHLX2o3/72PI4oTXkwNrM9afNfJvcqEQYu1/2vAg9dnMSCzsKivYfMc04X5g7+qSN
QGF2PvF5l5hYvVG+P5fSQD0tGmghAFk0S3NmkBqXEU2InstoHVL8RhaXOsjDLcV0LgsAsIvhcZmq
hsZ0QRa1Oe2nv/jisEknTKm0Uy3X9DqG0s8/lgOgGk26psT1WJFA4peJjcirvrxU9m+iNHvTKJaT
P7GEOu/aHOQwQg+nabNBMmdZI999K7Oto1tVp/uLCHCp8gF0sKInsBylXW8pXmVfQI3pkHj2Zzbl
a0apZE0LPbbacjJ8wuX4/5o48DK+Y2Dvm4LWizRzkcTSVX9VXiAsQPg1l2fiIVTULXJZLpKPHSGJ
mIH9EQ80KcD1ekSMQ6okH0n6lHycbXPgK1SXdrGE2J1BBgYZ9s7QUxOJ+geP3Q5fSEiTxn4cZ1py
HxiEIEfPtIERjp11Dllx361n+o6VCrh8ohkTGYt5QaLBsSHrXXny5GzBmr5qFcTS6qZDsq6/8JpO
24d+gugoiyr87q6AQnKnQU+M8CVSObESWi0ML7wliDaTEwtbartr/+tuJJYHsgOFEr9S1HSSdqme
u1ee+WaAaYwWtRww/070ULdriw3yzSrrc8bywEx6kfOyLTIgx2Ga4UXXmHQrJ385vUH0RIaXyrK0
xRLBLmAs6jAl6hIM/uMe1s0n97WzgsZ7CYKOGyjUIi1vokoZzLi0HcVaRCknAXarL3tZHBwUfw2T
NEyw2JNK2yPtq5BWY+67KrHec7ue4a/LlgpUE8vrofdSgWZTjbb7/IU98MPugeflc7ISjgiOV2VS
xPDA4tIKdpZZD9pJ38mmyYdkFYT0c66m7R0fG9+DxIrhlqRpsWXrWCN1X6qiKTeTBYIVtOz25cv1
D3PI+JN9bvuzYgc4TagVxCk2HENVage5cTv72NjDTDRj15Wd7U8rgX86pc0q4Fn4tvcvgA2QIUN+
xRgACxr3HT+zYJ9KFtw9G3EV4TZ15XzsN0tm8hRfWgYpurvIvQImRsKiWR0I6NZxmf1Qmzwuffl7
zrceMcPK3H+gZGNr8qiZWxggSuWUG0PPSt8ZZJPoc5lTPQwg8MfdLCImBRYLipUvcInYuxAG7mQ/
R0BlJDTYilP+fPLiMzirJ7G4jxScc682hz0iEbP8if1jRUqZD/dYN8ljIEsXsnSenPEP120cU54J
ZiSUg5Ogz4F3oe/DmoaufNlygVwCsZ8rf2mnMJaHaRfpNzPuGltxZxFS7OpqWQJBAq/U+09dLxcw
hksnrS3YP/jHmU3ju35STq4OioR1Zt9Qb34Pgf9pOj1Vs6RN+2lBc+f8fPuwMtP89yeLCQQ8SO9h
3GZMn4HhJ5wNfmtRVboXJ5PkG3L3+koNuW7AW3rQGV40vvQIxntPLUadnR5j2w1kdQxIEQm1npBa
40XkBtO+Z38H2pv5/M9yuw0YVXeyv9lzSwuVgYbTQhEjRXoYltcO+Wn2T5PCCc46W/leSGCpxy/Z
frhadySVR3XyJimtwBMvRIwcX0bMbrQxF3jcCzKjNsmyJAsxJy2klCR+jJePgza/IC8Zhb9bz8Pd
AaWYPWtuUvqKv/cWWjeAf9rKZp6VnFeG4XfqIA0Lo1eL7z1k+sZakhTE6AQtN1scR6SiB4pa1L5d
p2jKHlWv7400jxdY7kDUrR+fXlsc+oGwJHD79/O0nzQzOlhiui3jsAk+G+1K8Ma1eTbE9GIeAPti
noSo3RTEDICxmfkAZKSFz9oj4+JWtWtXNKRYejLpWWL0CVDbLVUiTixwNp0zuvvKQkCayZpU0iBM
0E2T614oBmkMEi+K8I5xCVa5ogJ2kdFLpKcEge/LuHezN2fWVu5/uzXqU9BdLy3WossXkx64YMZO
m5ypX05RbG1bUpX7V7VEEzuTta2nsPFUfD26ac4HhTeXH6BwUZZR0D/gx53CHqfMQygO2A42Tu+v
ANU1fgJfYneJv5vnn/MJgFGUXHLXIDeEg3ymJVx9tqPVAsvj42Gjdwt7NsfbZakJ7zzwAHwBGTHc
8oVSqmYaZTtmdXWQJ6Lce4oJaiYCO6upqSjIm+diM9cJgx7JMFltfljNTkLjDaGORzl5XMqEaGTW
cKoQFhKtQEJY5m3RNg9LLdqTS0CIaX75k37ABbvFM+BX/h9urP4UCzAZ4vWiRWyx9UAUCw5+L57W
Nn6fi9lb39N/vDGtCJqJBwygQaO/W2Bt7RO4/0M2z4bPmjQpeUqEhs3iExKUl3uDq61odPg7g7XU
pIuhRFKabnDLIehuzvZjs5XIyk8Q1qzF62rLFCd+hB2kNIInw3BFzM97Li6/UtX6ll+M96AcfAE7
5EROPB0GQH4L8CEaxunAj0oTJpz4QKycItheZZZsij/8vkAWcCXrfm5uAV6kpu9IDMykeXGb0vC2
/pm1GvkiybIs1+UWKwjqpZ0l9wdlWKiD60PHeyZU6fWMRY9+InKQNWGsovhI63pi/wqctr3SO2h8
si05egrwf8vr9lGBepm45XiNtVFrLH83IALraAmZJvuWSHXG/bE8NDuVT8UF6XbhPOJyGmsQ3d5z
E4eJ3MPBNz61ZegN9OZIQJu8E1fMHFGJcVC5QtEVaO8EAuX9RQSJZ5/G3ma3WD6H1NCEtO2ZmLpV
YM1bT/mxKyxtSxub0OhKUqZablc5SoQ2nMByPtpOSzZYwDiGXCjO5ilt1CYTDfhweZbRtrv6KrE1
rkW6j0r4ZkiwAb3rE8lws0qzUkmG+psp+/eNJIxHD+ylEYhf6b/tWc5Mp76xv0DYxkQNpjDNbRPa
TJoc3ctqnktPA/9SIidok4n5DeT/Zb9HuCezN24fEXVbGw2PlzEKbUdvHqwNRGhwDXasLnoV/1YS
NRVDLCWOw00/zR4izVYQFDfgK5pRXJ7DD0dx6KP9AxlkeIFpp8t1r+7Nj3gLgqzPXl0J1jRASpXk
jLs1ZUXkU8pPrHhsirITZSaEYN+Xr6vZfe5XEj0qDgWJwkt3uVS+5oKooWJsozMwLuhxEaPui/BZ
Cpgs5ij+vBxYslmCwn4jZpjRMKs/0P+W7wt2ylNHBrRCYcxuQpa/jSfyeOyImahGLVIkLbzkj7yQ
ia9z+ctlrmnN3y/pD3hXTTGOLRV5tTMqYYwMmC104RM5BkeFCHbD5PejcFtraKdLnAU+b0uL4gxx
DL7g+ydY0S0U3HppBrB23dkGAtl7H7eXw6MorofbCzjpRx6iBxbNa6RoXNEjD4Bf4JAkf8gVQzws
pjv/tpK4jVwU5lpY0q6ZxujalXtjZof830YgaxLIJlCL+MYmmhhNY63t+zNwp+9wJGsCHZTuTT9p
T+QLS4eUFurkBuUVXQXIS7tClNEoa6canrBvO8CIPag0a6sOH9lHSHVAtWAFkRs7ffV/3JJtcFBm
eMHMchbFJddmhMOj/8LQh6yz/rIHFuIIrxR1hO0jTZ8wLx3FSR0/M2Gt+5NiyKN/bM3kJE5zjwhR
307/itsz4ESV2RLdM+sSyidEcaEA+VXxLj5aS1mKehbkk1v2pi3jBd+M9I9lQ5GAFMV8RazsW5mK
I5/DqoJOniGFiY29XgsDGOBdks5irlgW1egfu0RYz8EjBSLYnGnGckiZ75pWZLJfo5Wf1kniTCTK
mZ/g9P01oHnsZhQS/6Z4G+G+e4MkKgvSrxYY0bn0YZgQgKKoBUkMhpt7yn8647CgRDtQkckSJF1H
a4Qb4BhkivWlM5uT2ypQkUbPEUmaIy7CAUmZMKrIN0ocZz22Ct33PJQiq8yjpan5+IngRH8Ie7O0
tF5Lx5VTVqHiph/tBWP69wii4wUvNky/6D0bDjP6Jej1dRso37oOarae/4WSgjO3HRDVf6ktP8Q3
24ChLXmGEltlEJ7xUZvsrNSE0CuhDlXSMw42i2dlLJzqqcAo8IzPPafrTNgl/r4Tjwplw+N1CUYm
wWuIVYWIEucFr0OAcS4HDPdhCU23rrDzQyDdRBFLHEYCg9iWZMTQIe8F5uVngA8KLBATQv3Jg0HO
6kjD9mO6o9os2v8PURqokBe1QU0xxmSsJaC0C4dpU8BpWarPLHbTOKMe/p1dNwuXKLztuVC+LRGx
lni2UM4Tc1CU8P2sy/4cvi5Ph1liO+/aM1Yb5k30UrJiaceQOeyp0vpjOD54GGAI1iWb/e8aApHB
LXsJJCReOJq/NcWh8fKi1tE2QyoZ0mb3JqRyfmBzwYqnhA6AZe1Y5CI4cnUGQo3aCzpwroyRbnlD
xUKJn6Mz+mDs1+6VFAicled6CSHezlLtHvL+vsWRGTk97l3cZgKrxveY8FsExP+vyi2IosNgQcys
Bi0gs1gR01Lq96WmPMYsWP7WavvPXMGrQ12NIrgQe/KjFIoByKRPhdPUwNRP4w6kL/PbVDXR+fBG
sP3rZPVJQe+aT11SCRq9HekFJ0iLT6DpjvzzxTh4v5TYWbaxTYuRC/r5lRuXCNEHC7Xak1zEZTrf
z6wlghl8xbsxLCiStIgjOUlvuTDQ4LFWKXTmzp2PvUTgSRqEBBLeddu6bdzDIdfE3s6g3QK3Ngoc
pjN71zetxfUAg8PAwJrh2z7uTLRFR+kWJJJxZPVMnLnb1/MxAgK4fjH8qauHWYEQ9v+Opu7q2E98
21oMjf4Upm8BsefJrSw9jjpdwBoYS68mhnWZPQdL77b/FB5xYr7vsdFCtXkQQnUAukPBdt+zNbdi
OEjEDXn8Xs/FP1E7Km9kxm9pJEuTwWqOT5PTepoy5MbxN96b+GA7BS4/VBWVhP1JorYVQHE2ojue
hzOHMQpbCDrkk2hHTChY0Zb2e0+r/CQYv5LoqAZAsLBNuL/YJv092JYYDeuP6Yoji3YzBt9Oh7+P
HRnvWZtgPxbPsl83gojZgqrTjjB6JyDR19BWYyVnAdy4/ApjJ/jJIOVA8dEM0tyIkd+3urku0yIL
jBSK9npEVCwQO+yUoz3t05/YxWDeeR4DLNrjzFZYQfVh/3NcYbDXgPk5esxBHDTMASfaMK8tV4+x
LJLIcoLDCwA0RAOAu+X7DCWiaJeH4vOa9GFRPg2QWSsvE44FGjlqtWdWOLpCOo7USFTf7NCH5dw+
bj6f96qzAkTp+gIjWVO+bR9y3wRbeUe2XXv32cr+1f36DmnBIe0mnPpg+SvAYM06VRNrLfG7bOpK
/0DB8C9QyKkd+YJ1g0tReEWgkBZ4DWaOKdfZ6DpGmGQoBYoROZ464urEIdbMs3Fcr7NxNl58Mfhj
R7YqXAPp7EcR721/qmUQTWpbAVZRQSmgY811vCLwDsNZ9qyV/Ogl7yZsERZ58Zs6CJWE5QtLzupW
X0s56MVOhZyDnPCExSt1WKwCZwRXSz1/2vAzUAv+3PEWy+o5vypZ8PiNr+Xm9HoOiFsuGo9EOPzN
zj7xqk2KzFpI+z449kjqbfA3z2nfHQrIdsLjqUmpQRDnLgSbg46AQiQjuv/BnwVULIDIqRn+Uc50
udV4RQIeN/2ZDPR+bmSQEte6SLEO9AobxnVvMysATpmKmhzl0qsWLOSwOyvDnqjTKNsBLNTMonK6
mxI0SX3rxc/XgS6mf78cAY5e2BKmQGKFtgb1PIgfdZGxJtBU9ffCZSeWMCjUGa0wZ3GVN1EiLanY
XEmlOPiPi2mtz8uZK9Vi1ueqo2/jxC+lV+HS9yylERtMrZKpx82oA5UOBa7Dmpv5qv8ckvxmBYkX
skFL36lhLzxDJu+CwtYfdCLQZwntSxQ6qks+qPZr2iHyCfghyXNbw+ac7I6DNdyDec1fCX/ENr9J
znhOprIznxrqAPPn0w5FScQGeE8opbQk2Fvokt5z5yqxfyCrBkBNnwolCbmHN7mx4DbQ2E0KEazZ
KopVXiOuRVcUhfIS0/Jm5I09hDUWh9UU5UjEGUKxqQqBSYZNSs7ne8VZVWs2SIjVa/KmN2FTD+8F
cynTIT17w+55LwEQ5sTtmOCg1+k7q7FVdLEhc5y00SZsXwvl60KPhNJaHxuXj4E9TMpNF848P8ri
vsuAdUJXuBFqPmVnVxH3JDaJYSwDT73bFIQkyzKr8Zg9NBMg3psjGPwX1Q1QcgU6fckzA4HO9jtX
wCjCgDuEvnNAbgn0Xjbyh0VlTSGcNxjN+SYuZtjxk8SqICDAfZqWRIk2v74uc1sjZuobVDVj7olc
KR6Z2GXL7jjzie89IUvE2jGx2IkiIzs8wvu7ZRxICgKKvQ3TEPSbWAtoVc5SjYGFt2Wbse3g9hNQ
Whi8EoiJ4eRrB2CFifAwN4zcNE16JvtH7tBiOoUgkGLf/d7ruAXCgmf8Ht1AuiUTh8QPLwzX58vh
hzu58EC8qGK64jkS/b/2TbTe/5hzAaIC4M0bDAW02mbth76qsM/K+4jE2qHjwrSD97/qlTCg+rXu
JwwCZp9lIIU/DgMTbnYG9w0Iid3uaBCsNM1oLLieHSK76ltifQHWNwwcQtH20KHruCQ6p4PZ8AYh
TcP7wXIzVALNRcJvG8JYTvTbM27mhndh4lkc9BtDzFVoK1DH6UQLjlfGPn/uw+r72sM0NStKCf+c
0Ij2Q/IrrOQNV56xt+Y97JtACVSoGbibiOiA3sPNrvQpad78FsbPjQ/a7iSBxtYVWqdfYCHtAqb2
z38HgpjAAX4x/Yup5FpZmMmHft31r62iYmCGnmt3PVXief84mU5DjgNRnEg3qR2o6AFqrng2XUPW
GPJIaNzrPq9GYP6FVFqVfB8tfL1NVcHcY6JIPN6KOsXwoqZ0yqSPu8AzeGaV4yz4Kf34FMxoz+1U
XDOfzJiq2kLow006ACeiNkbVlm5QmhlgjvwrQV7THjVSgm6LtKILUSzgChaNlFqlf+OG/uhje8NO
iu5ASTkAXDn2u0BrHGFxNtnOOHtP7JlcsA1MOaEJBAwkwh1YJ/bq8gy21feZmYYK1MRKaJcDyGlt
+VLOEzz3DbPVrC8kyRMPikj77lIeHc5f6yNVe5pvrtX3xjf3XXeGOf5CAU50OKl2PO98ki5+Z3b0
EDXbRg9JK1ke/x69Y9k6BBSAQVKmuV7QIDzgDIICYRhqnbBngIJAC2s5s/ITpYgiCD3z1zs36nzq
D8LIx9kh+lu1kvxVAiwerPn2iLPheCYukZhcRkLc3DvRPhVpe3OJzUbDEamuAuN15dZpl5YkZz70
SJ2xauQTzXsLUzD6ec0lKThZO2OiuXE6Xgv0MYVmhHMqHr7vN0WeVmoxxg0C5wGGn1JtXqR45wsM
m1BRjgKeuIuNoXcxbvXHipY6v7DX8T+xFJnaHGXZziEjDAzG7iUPp5JedILz5do/d8dzsRcUcUxP
Nzh3AFuZDLfn3awELTGyoZZYzBgrRM6If3hXTJ+wWqeiorqMKZu4tWTttA7Gxp5/BRJg7N2aTftR
YnxoRR5VDJYr5CoMoeiAr0NrXOh3rQ7kk+2rzTGxxhBJ0VplVeUaa7i5jc29OKPVIO5vBM3U2f0x
Nq/EeqEdRLoAzRGXYWOoMoWbtdBHW9cUA05kXBPlOIDAMQZ/VoxLOkPPh9DWjqouZFUm0U772m+c
zvBd+eASJSGjhU5l5D8l6tYvKElFMq+fyUT+o0vmj9kF4MMWaN7Ku1xFW8tXB4pQXiSb7zxWPq+a
OUzAEwb6/cZ6wNXdAHBx0p9hNPY8AFEMEhLy78z7xsj7WASBu1qbY2eNBd8z9Fcxjo7db2bfqkow
Q2Wuzmg4EZQ1PSFtyXomcVYtXIytUn28JNVj1NGQHDUIqOEXMtlQuOLq0e6ouYweYJNRD5Uo0nL9
3xrzdc0IPNtwHHoQ9heJoeTYNXrGRrs0uKUJBeTgdbKijOKBaJs3cc5lv3TRWanblh3wzd3d+p7z
a9FCVDcVfWEoOvuyxa9jIH6OPiO/19zYAJJs9u5KBW6/dC5T2GBHF9hYI187sVOwaDlreG4HxjCW
ZaP8T/BmcnCmEZMwqO0jM1H1cbUKMnjzjNUEWADyNZASunNzUYTv5aXinkHbk4x4bG3kIWlAR49r
BsG6t6ufFnEtDZpMj9miD5+Q6rmfYXGyBz/0N4rJDYmxrjdR/Fd8gZC1CBWni45gRo9aNSoqhSo8
eCc4sZPB+NWVcsKSDBdMCp0iG41NoV/uUVsf8LPplf6WZGc5qT8R/QkvvZymc+eEqbQhtHla5UUt
M3VmnpztSMNEisO8HdajQ2gvUfaH53VA2WqdCuSuPoxklgjimqiu5WS3hmsXj/3Y2t6U2QcbFs0Z
AtMxNc/dYqIkcut4npvRLU/RsvLJndgLipDM0EhKm9hyOobSzHhQ1eCWamWM4hVzIKMtwCi94a+k
D4bpVmb8X0fBa7jB7NcIosxDxSwpKj0TdWKaGPo9+tIf5dHeJ7fcxLnQSdr4hGE/bIjkD6JloCfk
LmhWiV8h0BOH90YmtplkuTdpN8RnJ+hIsWdMfriV8W6EJjUv0kqJYKccBlMIHULZoBPuyMTSIgc/
3Z5ejNOpWWpf+ZkMwzwHKQ02XVsbb6b+EEZven8sRBUHOCCzd2F9+VwlB7B1BeuRbh4qjRSrJ9he
RlotJ0MNbDnsc3Hl5eKzGowpxs+l9bVZu/DgPErXAffXa/IaKFWUtFOR27e8orpUQA4DFHv9kKs8
Wx2XlDDtgwZtIGxWJGw72E/jeptDCjMntEDOljG4ES8LvBRv/+oDio0Xgg6UZ6I0puhjilvMGMEq
BWxOt9lP3lwd+har1QH1W78MAGgyZ/HbZz30/24VQjSLPPdKpiSQ6AAJ2hMpiD1IgDQjqET1FNp3
XIijnFDPohzrxDHtrITnwEnGn2OL84ZUjfBg0lb0Dotb9HhQZ5BbPLdSuAZjlJ38+i2lv1J8HE8c
JeqC15hAkaurfxr9xqt6p5+stjinJeUrEHfMaF4ew5x1C/vuhvwEteFO9iVv+BO79eaRBzY5s8cS
aa0TjSEo1b3un+qWrwl7tz6GuIz2CEg1MMl4dPHWSixhfX0Rf9kqacHzmbIdX1aXPBLAdhebEWsE
q+e3qY3FVJHpeqc8LsdGptMKufz8Or3K8VYNrj2HbxAgHyMczEy2ZJQ+ksF3SS6XjX3HGQWYyeGl
Fia0MPOrfqaJu6J/q3YhSupcY8hKumjrkF1kqk3cELbN1E8IZHvymg20p3SUhoPzGcXoG0gCEDPt
p+/bv7JV+g1BOhMc1MVrlUt2hNhUurYONVnfdWlTZ8GrDtRME5ZdKT6y0nBtV/FRgeYnUyQ2JV5m
08boTYfK5ZSd9eT/+B2YOJfgAHxIf+4MZ8+rdh9+4k2KMCDKY2xI8Gp5pLSieoMzhseA+Im1JoA9
pE8uteVczOZ2QLRrSSaQr1u8tjb5GB17Ir09GoWcHnbD8DHLwIe1mGWXN5bZLTlHab8nHl3LgOpF
7T3caeDaOpyRWGoHlc/kVW3Z/zdaI4mGqwID1E0r5xpws68ZHbNkPNs9z4lbSLUOPRFdrMcuO0da
7X//mBdD7L34j8uqqbuepbTNaUkiPet+4/RAkNrjD/qwsWy0czsJb/B22HZpe8+PgpBAw9CQAKJe
D/intLkRkKXF66EYfQxEK523rYo1p/rJVRcxKCRAyhtMKzVp4+ZeRaIlbsQGjxWqZflOFoDAEhv8
ckGR9XzN1x1rRoe4QA2xCP/uMeH+/sl+ZMVOmzZB/PnDQNYdZeMNjLuB/j/ZRUMFljYuPBSr/tg5
L2omUNGQJKtt+1lqpZzBNgLLhpCTh1p5YmZ6kKKDSVV3twIxNkHhD0bAi/1hNRCRGzhOKRBX/dU3
SGabPhPya67RVkBETpa4T5U4gT2oQ+6G68nRXbRF5UX6riMlK6Bv/nGgx2wdFfPaylHWiNVWwC//
pF5ddfXoszg0PQquqfa3GmpSa2oNPbUN8U93t7nFKXO8aQLtGA/UdIGbelfmARsW2kN9ZO0okEdL
5prCd9u3sAbQvxn2I+xOKCT31hnjrzxVkJbTFymsWNOIvf8Cb5hn6YJE/gDNr9ofBE4h9zbEIOZy
CgsFWUM7hhenHr5ztZBUV20md7ERVkfINtYfVm2C8fWoi0hewVKHsxKfzUyTQiisX7SCJNoar+nl
CneXFFTW9X6gjgVpoJou1ONsvUqiPK6+2nitTCbLmCBkrV4Rg8/YbBC5NbQsId4gz/jI23ppGr8n
nUVgOztnjdPB8JMWI9iR46z2DQhklggbIz1LCqG/oeVrlwreugT/VIsBmOJP04PualfGJwCxxAit
6PcXNxz2LqyG4I+zI2z5k8s/UqUtHxr2+PSGKz2FI7HirI4K3TmjsjQR7/c/WsBb9WuXHOWF1PNS
rGaR3Jkwx7LRP2FTh+hBILQZK8eaFaE8OZ2CjtQZ43Nk2DxXNX18wTf7IZsE32Rs1GwM3CWT2WZh
5/SNeYGhV+7RNzVXGohow1XlRbiq9b51tYRQObeGO/7xgV0C6WsdgSv229nUfXtsgAmg41J8V64m
gr/dRl47rl2V2xJ9D0UItQwwgWXkbrHN5pIyZoXKQBMTAEAcdYE2p8H7aio+NSkzLPq4GcdXyXjF
VzhN+MwjqQFjNtsy3p+csw+0gKwXpmYnuNxvC5Thzsai7Liw2aTEe5l/qpwwYeAU09+UM6pFDxO7
2iIXJmB6Xh78za0sJXZN88gtbpkwykxTrHhuP5ARo2eZI8AP4MKODRMAjQ5H2ovXraM/roAGZzJ9
97tetMlZC9/Mshl3UqMtuTkSV4xeemG4QUyoSx3tHvJ4QUkZuntYqOlO7h+wyFmNxOyScUIcokuG
5WWE7PcxGYHGDD3XT0d4Aywpxyx883MW3TNilOAlIi7VzQXZX8sxE1oOo/TrJ1/eyZcwWxf580MT
gH3YLMKRWl8Lo+OWG6dOs3Hf9nbQPWn0JUYa65G+9vBNMmkYNQmWpzBsv6rDwJn29wK16rU8EZ1C
F8a+yg4jG4HHtnA+vv5exmcKc63hRDzAJLLEXk8DCWFD6gtCBzWp/fQjuvF15HF6407/+VhT5Kb7
5tVg2ILjo14Yuowvwd1tdABqp1EVdnyN3MJSc4YgKu1BplV9u4F64hgrYUpgm1cOmu6jFbNerBNQ
0PO3oqrwBXRkl7qRrO4tScUQ6SWxrlL1wNU4eHOs+MgwSPybwzhlaNKzEniuAnir8gCTfJw76dyC
3CrBU26MKbzPqQhQH5rnWfqCzWcZ7BOBF8q5qvoV5jF4E0DeHoCRaJmXTvc863m6/1W+7VUgf+N/
ULFud/jl09Sqyapb1YGhhbvuDQlbYxhOKkrA3sUVLl4tIwB5DdimMfgo08Ro90OMI8QhCQsMzAkb
R7X+rQxNoiQIrolTKuw3HvFWjU55oYD+HDEsLpqp6ZwjwSRMFivdx7CCDBacqG5wGeZAmTZ7w/OH
y6Og85HmxDa3AzjBTaMnUBqPCEJtDqCKDuLi3AoxUwpmo9Wc8784WiKJNc/rBFpdBL83BsePKylL
ZXx/leFycg+EH6AiDgfiCdTKLBGkMupIeuyZBNTpH72/IY13Y5JT7THSrrNfqxfY1BtpTqVvcMXF
GKDDDX+thtRQG6eaIIZVFDFU8PQVfDft4pyn0WcZqH/AfUnvNSjluNMRK2e+bAhe+DaaE2LSvUnF
U4YTwXSKg3CNXJ0ne+Y63uX9hluhJjWNsHJQaWv0SAdD9G0jmlD/4SAf6x08MJQ+ElxCov2bn2sJ
bpVOqurtmWhKEvTQv9LzprSm8OAqRBEqbMrOXu8Vfc9typYBjQCcnQZFmp7oI1h+AUtxiKeRYu2q
j4ztJqihweAWowvnoOhDDT35tu3A4fi9S0cOfoq7zTldsjIfOsohgPCmn2sH6jXxG8+V+lVHihRv
+g+py3aYQi9MP46ndVQojScLfCkAnX4N95Zm4LYKJ1SUI6EjWYcZJ8eX02OIlXeKFjIlU44xLwD3
BBtE9Whzc5bf1tD0+/dknzcRNRaY7yZML1swgQLub7BJqZ0OdwpPjPsSAuFkD0C27ChDStmsgG4y
Bg62BEB4mYkDAzXGMX1Ft5gJ06a8z4XV3J0YZla7p98WAyyu2TRv7R0Q2qKsheHD8bwbIjnDywXM
BBoFpNAjEVv0Lk1VLyr6I346m6WdcXyn0Z4UkufmO9EuUNgrq3yYQIzTAK+Q68s6BnsvgtVmrcUU
25pOUIDfoBds4HjyZretoTVLYjtyXWbsqrB4My1CsQwXw4GlGHODj2P0j+ZNQTT6Rx5PZW72siay
qRKBgRyl2/g1azXsgybCz1isqEYqwQLNOO93ASplSQRWt8N0VMhS6VMlFOp3lqYm6S5RBGK2HiHn
8ggDh5TPRbIKtUtDmcPaZwHP8yJ8nKSPjjK0f1vJZ2CeDq44sEO28gUFk+bYqeVs4ri96fTVKQss
hNVjizMKiqbf37gAs6e4cdIHbbUejJqqnXTfqBpDy8FYsLai+rVQ4TmST6GNlSGhU29Jliopt9XR
PdViI0udotXXXpRZfZ4+xy+CAM1d8na3K557+h0mdi+cry8T+3FsaGqwm2rfnr9asibIYwL9WekP
hh7xeN3VZwoelYst2BSvEmoL6H5MMflR9Z01OPR0lfqXIlwjoEieljmDAaVcaZQrbV7OyXjYLOot
t8F1PU7V19LgQXm1V0DvIUkQZSbzX5adMfZCEAmuDNZE13WW59LyPzyLAihQEbsATsF+AhPcZVXK
Y7SOUmQQY/Cr3Q1t9Io4frsltDi9GAILpxVYkRWY1ijf4RCRn/3AjX6aJ1DO/ofAHKZdKRPnIB8l
Os5/UyslcXXsKGMKsyr6PduqfZ0shgbTuG+oND0FFo+OyBNhJDqFu1ierJXpsk4/ikDxX8u8FNN5
qhn1wLyASqvG6hdESTe9r7ayt/yyp45KX2YCSvzUoHO/JKZrqNM1e7/QetWMADEiKuMGQpalLXcG
Faaw1MUbtprsJINBzh4Q2oL+qDSY6bMi9JttKxMyhIb5VLeSdRVML58koiKNJg+u9PH3NzFhCzs5
NtriI00vJgQcpquB2cuEFJe4rnWpf0Qwyl5IrqshaO80SNasRB71uB5tc/eBcjqb9TK9uyiDjMOH
gOuqOVFNrn9IQYRfPPdNWJg85gKj8a5SR1zrvZzBgrib7kYOpQM/1UcZSPTZEgEiZU2kmHQwhtkG
CDGrzWspL143ip3Vy+Zebau5lbNqCn5UEPC+RD6JrhXIzoUX6TYS7XMwb5dddF2HdvjssIhQTw3Z
xNuFcrDvt6O6h/aTfEGVb5OC9sZFOT2YV3OTsGbgGI6EFMatizXlywpjRQcjGqMsqLcGxonx7q2A
PHyylq5CQlTYetf6jVoRqz4xAWrBY9UjNZJwnGG02dIs+VjvYj9qV01FV0m3pQxfq0+zZ3EbgfzJ
kaKvFLS4UqNZy7t67sajZ8eQJ9Xkkc4p54XbRWpHbg4Rb3optZPTBU4+q+gn2xFcTJCLEOJ1MBJt
rZ1lNNuMksk9H19WgOl9Bfy4Fib9RZrwzOWDOEozzPK4vzBeFOAjtP3eX43ckZFPUUcaQH2pyJ6f
M4SXcPC4oU9+s0BD16JjmAoJq4w9vMap0zLU8Pu7y/RpAPIVX+1TALJhCfh4fi6rdars8fSY/esc
X5VFdRy9g2WCRcI8p9UKy5ze5BpDSokNT4PZEPOZhQVbBesKK1r7CXa9WI53p788QPZQYNLtkBzz
I2pjI0hRNtDzDnXZQfLV6PrcQ2ADkwv7880h7+wgLkzXN+1ItQChO9q2R62hg4fp69wh1pFF07V5
K3GbfualVnAHC/piRRXovD1L1BGIvKHBRgh9npLMahvSf13gYGJRbAxqM1FKkkJyNp57CksPCzl2
APeCo+RiRRuP4kXfRkm5WfH2Dr/kjw/NVAg1/uWaeZJk9dtpgx62AAB/uwEDtBcpQKy3YAhmzPRJ
CEEstXt90IS8MAy1NWcGeKOzFU6ilOUvzlvEfVYQi/3J5/v/u9H0CogpkfgcE15PBAL7SBauXLL7
fo4Dsk8sIwPZ5QL5jS6q4OzNdF5ixVjSS0L7yXUMM86DuXGs/9T5sNUWym2jGWAY9T/9nnvymwcu
CVmvz1HMgU7oOz8Wkjinw27WweYTaEB02wpjgj/BoIMakCKwi8niTPA/bhLl1sR4FB9jRZGcFLuB
X+XaE7Wrw1D+M8udfpL6y7L+c8MMcZSXHkPzBatw6cpOs42PAe6vArCu8fuH4P2vxl8+UJeEPk/Q
icVq1PK+U5tVWKeELRCwn4XKqYffkYOyXDuLCLL/0htWk7mrpJTClfbRdPRJ4slHzb0t6ZJTWEP2
kTXTiEfp1mcjmqjsNOt1Aa2oDWLw3/4RdIPBBAspQOko2kEFrdiU4TtHUq99U+WRizT13Q8PGRLL
ZsInhLJemWHOSnWA1H3+2neyWFaQWvDCwyCFITKcmS8VavG2O7dx9Klqyhhl8vKUsmnqjKg6tdkq
ABuflyOf4sFJwtI6TJJXJXGypP2h5v2oVLnivE4SQLTJtLfUbXERdwe3LWioFpPDpqm6h4PYoucn
LYje7F1OfowDycx6s8hon+4otaY0tNcw2dO+dMDgDBJZmD6kVzcmi4bLOEb2gxkeZAHuoMFXDhI+
qa94eRnxHPtKkITtLGGXtZtAwk8TlU4tCENR7+YOTL6+zFAxT4gzpJX27yIhHx1MHjPrKzpGC/sa
50U/kvYAE4e2lfIP2QCok89tLCMO3SkWkOP6N8kL+imoSHPH6SfFZ3F9Op0LITVQyBUNT4pTJCXW
xON11dhcODznUM/6nmnsZhux72izwsMmHRICFEENaW/ant8JNUm9L+tzhsKuJmxch8WAGz8Kp96C
sGcr/H2ipOuNMeQN9876AMh9HmL7P1c2wBiQC7DLPKV+OhuRLE1N0cYYZlKZqUS0rxjdR81IoG9k
TIhAPt3jDremJcWYQf2qsGWWAxFHP2t8RIU+RDt2DHeAH0hFwXfka1pE911DwAtuuyolC0tJiqOs
KxsKuEPDQspza6Q5J2rWbRmlwMDpf71FaHbR0pzb969Ojn180cdhl0bpcd4X2j4XoCxAeG50qMHI
bGLTAbJxfFPiSMwj3T4aHXvPxTQvD4XdFsxUAslB7oe2tsyQX6m0NiK+gA0l2HJWOfrdIfGiC8t0
6T542Lyti7GtDFDbwV58gsU1PcOcKnVUzlOeBZ98lNba1R+uKIPbHM6q3RcHvFXpLiNFpHbygM2Z
ksJZs3HgvA7VqjwMtCtGr7m5wBax0iI6nBXEFosy9vPIA2rbzcLNw+m+Ypdo4rl603bi1VuYjWKD
s0PTJdXiB+nE2QPdMO4PPwgfsvCm7tYDiSHh6/U+83lJa194KwEJOzPo1qprRG+5Enim17eIMXnN
VK1G0CxaiZcnQfLA4hxtHtNGOTi9zk+iEJ0DxGil3iZ/lvFHLWVzav6mtT1l/GCeNuq+WLb94j27
4THX59N/FlShB3WNDl2S46v2tF9FhbMpBkofjRWmddAyRMDKQ4SeurhB0EyPmBsnZ1j02Zn63P36
bSjofYalK+uoIoNY3waued2f39Tw99Nk6Myn+UZt/mTUHDyl5ncYqn+X3oOPEvqO6EENe80Uc7Tc
W2c8w4Or56AmDFWVjyS+zfczIjJi/WMiCHo2CNIeVuJWmASJONvzyBOTsQ9A/+D6OIxzn/gitRJk
63plEJXSLJ7oZYguNCQgsp7jWYSOkEMgEqvDRpofqgtI1QL8qOb7JnaLuVP9BQ7RxRI2xAvByiVA
dWpsDsqH4vZvcbrvi/PosUdaEF1FTrv9dQhMUmtCyP8CztbMHbWLp+o+bkW91G1bOBVn2MLsX0KM
lBtWca0M5owXE/V+dM1kLa75X67op7ZsQYGoJncn2Gug3P1c4cZAKxQRnYABX9pV3AtBtEs5UxLr
FqbARF5jY0/Bu0EqPmGpUQiEgP4LC1zU661wz3ZoP4LT+/xwgxYU6WXQvbY5z5UKLmwT8dRZcR09
MNEEXrQAD8GCam/NGZrvhfkRisTHtUMeBZjk3Db1/7NodnYN/kOZws6IMB7BMYMsIF5/zidAVsGm
e2DnHrLQuR7yL5hA+WxLnqYR2N2Aa18HwmPQwGIhAzlJkixQz3le/7FMWZhOFS13fj41hxbpW7DR
30XH8bo++qSLjkb7tSqNXFegwZdGIvHyoiedHIIBFLkN59w1Y24QcxBPcI2VHm16g5aksO7SKb6U
gZAY5MI/Ky7HuWS5OBnQNsZjmYKTXWIQjb91kEH7MDAHCrhM/PrvbRTpN5321cg8XApDYWY4hSMk
pZn2FEtJBgwWnXshxvjKEYoSo+aVHHseD5Ed7gJugVUTGmVLKn9398wcryjRLWmMNa99lNbb3xS0
TGPNZwAIIaJMqNjK+1Jhw16KJ/ciOxd81DG1amdfskCG40DWy1uZ07zVYeBWADEZFbkkxJr38ttt
mhft0jeMBL6Elti9VXZNfRxSaZVhe1XDUpSR9c9aUHQja1bNFcCg89G/JH0P2ZWNEhkqfHy7zM2/
xO29s9/oenFSD723wmcFdmcdncg3OJMLw79KKFdaGFpVdfiUrIpqXb2GwuANYiNCyOyGmP5FrXtA
HGnrVfMfWatEW4S9WFfUcBgd/c72oltyG0BLV9YykcX96dqJk2erSO+yg9ArQsTto5GE/MiV1SP4
30AbHuq3N9xPCixE5NmITIL98bceMeKC52F9R5EB8vVhsBF/bE0SnXyBSlxKc8WV4E0ysOig+wa8
Sv68f7ZrrnBPRgEVZzboYACC9Ac++2Syr96YcRESN6wcaooDI/pQk5712fUu9eXOaEfRTSV/T3A6
6UXLzUECaEtIxsjzcJEHfn4v5jbZhn1w3yn1K8H91ayAwgcdJGsqv5CPUC/4w7DAbR4AEMvvKhj4
cb/oahGrqDTT1QAkVn+aLVxzyiagPlrKK6BP9YWI61Jtab5dkzbScnILjlx8q2LYC8B4Az5e22ci
r73PvwX/BsNdNHwCBvWX8vSTIlk/qQAOi0IhHxKxyEu8OeU/fo0MBFwvyZVW5iuJMIxbCjgUI2er
r6r0MjyEE787puO8H35CdxtSTmAfung4vkcLsGt6K6ZZf/qNJxR+oBislS0v3ZkWD1h+ewGilieV
zkoe4LDdnKzdNW3Uwogm9cGVCGE+Tlg8RadNaoqBIDGrAvJ7DJ08GjUYNdpF9yMhK7GNIrICVOe2
wwkX5rwhHJO1cADXMaXCjgIZMA25nwC8UgQHOdyqEQrNvuM0+mnJe8acKFQRojfHnjby8WX/+M32
Q+qvCU+OoDRSCfTjcgFkEwaAD+LmF2oAt+s8S0TqqZa0n4GgM5NDPM7pJqt+o3LHytHGE2YnQhSn
W0TEGn/DkaK60njb8fX/566ObOHZy4Jj6bcKh7YN8W0Sc6/rXkCPH/azG6RL7ypNf2b+rdrACQhi
+1Xkm+OotmQqMDeFmy1sOCNFTo+bACWniebfZp8XMqt+PrIjyN9tNZkWOE5P8se/J1wGJJ16C9TG
0tv9rhQKO1zOQsjdBhaP7Jvd6+WI1oyrFJMa7u1Ab9zeThYt4OqAjGd1vyxILj0nsbNGtEcuh8N9
ROutvqrt5Vqn1XNYCXRCyEFNmQdKwyfOaFT2wQCa+/JMV1RpMFWH9J+Yy+GrLUt1DdjNaHnVvZUf
5U8+tMfMj3ArmfI8fVTVOTrVlFjqvfvkLhGvj2nFufiNiWv1iRmdIODa38VB3bgc0hMRnqQc6LoY
Pdo1dOi9gBUGZNJXaadXCWk5+EI3fEvHxzup35RestP92AG0AFgq6way8bia0ZUYr2NGNy040PXr
xDpNUr+UIIkeSPFfbiG3TN72LsYlhZsT5RynBQG6HjTRhg0FMTFymCmz1I28J4pXiOL1j0EI17eL
wnnP7N2XocmpTEImWwZVrWZf+0XgijoYF6iIo+sPwfaBfeHkD5xj3t6AlafbM0oh1GdRk2H6Rbfl
HflDW6JLZbvZc+LpNqyKY/VGcbauw7y65jpYDeBbMhzpmQhOgG+6+FeYr+dR/U5y2g+xEkNTio3O
qd61coUWuymyjLzHccI2vfx20VaFGACyIEqPjyw53glElzhPSooavmsZumlOeCkK3anqg8FjaipF
K0huhJZ2GX8yqK78pPWLBth2dLzk/BlMHs1O9RqMg0Fx8LUQxH73tQCYLLkLp3vv5RHmRzgTTHxB
LPYxs0WOQd25ylsST5Gjvrb+IQJhWATvJvLPA6kCdJ9ohXuPy4qJRwW1qqbp/g3ODfxl7z2eFgdO
EQw5++LPiKJVJKaWJisJEVSoAE3B4lyulCZIOQYLOzSLZVce0c7AU68ezZ6e5DAp4bRzs8iDzTRz
8TkyjQrQqiLabKoLJ8rQltksfjSrixaOXg7jNTB+0OREvYXijSJzjRwhq6M/Z7yd6uV+7ZhhJndM
IQZy6WAukoRo1sfpHfXG5dLv/LQdMW2Yp5/qySZ/HMnc5vr8E/5IHsJCrxwn4ffGJddWWIv8XmB6
fRztAt2Ol8cNFs6gDdDtk7An4xaW1Iy2cmLjgrKYt9kLQKXTzHiCC2jxphhAYjJ9TM1EdKUcM8JX
UoRNJhFJtlrDASnUrOteiWCDKGKlBaL9bDKURTlAr2vM+CwcPWFY6xERJAw1Dd8xYp0yeGEFoQb1
SzMQ02l6/9jYho2K9vuZyi4jK3PWs+Tf96qjSJzl44DGOVYfUQA9vbhSPVZu3u8knGuQ0UekPPOO
SR5+nur7BUPEL4l+GEfffOrm07obxZEmMnlB/hrk5Q5ylyHpby1EO9ZlOEq5j+L+QqrH28khnj4/
hB7Bnt5qzXSTyDGELD12ZZM6Eb10ZxFTDYFZiv7nQos6wwfBbCH8w70yg0OY9SnFGwZrRuKlkWeE
kkku8adN2PfMfJquTyxGNMfDRD6lBE6cxiNgefmMDiUcsXaCvWPe/BTqzvc8AwHuVSFsAaABR8OD
ldptqlFqAtAalOqvjGGbmosSIFUKCRz4N/DN92vEtuB1huCl9tPfyAlFvs0Lmld4hAQzENw6c7ef
a+Zh3/ma61swpKPiKbs+mxmVWWfwrnO2qSYHZGZ9iCqWcsmZ42S9aYP/StfkNGG6PYKTup75ONFR
bCR8z5GdXdNfHcjUT+wK+GUx0zxnBTTo4lQvc55eps4N0pjZPXEkMw0OPNZdjht8LjYJjdA6R91u
slDvhMlE2XnSxBOUFpfpdGfERRooETAEQV7kXCBaqJtZXrhc/8Mm+O38Qadwx4qPSrprqU6jeSg7
erp0CtnVRRtMOkpBzq6T8JpHgQme1vanezLDAiC3YhJFF2VTF5tN3tCyFIr9eNBXQcRw/s+jsftP
TEwf7AnhHBxpoNb2KyagFLJ4mEQV6h8KgKyu3sq2I4+SvQZIKcU2lKd7TMbQt5PK25nl4+qb/Q2z
Fq/KN+t9b6f3t/e+ENJ/Wb4fFw1f+7ORyUSUFoAiJpKyRNs+Tb899wz3rJWyRxCdmp8J9GNcDsLO
gX43J9+OxQUeQkTlXckX+YkLKiXNH5240rhB5H9v9NiaVxtaN9c/QcpCC9cbV3R0vE8YYjLbDhtg
Q//L6htFtJElcXlmfxFnlfF5G38qbEifEOVw4XkHmg0TxrVAstviHTEJqSSv9+GxyT0k7w0Y4xZO
yVTAV9QHABgz2mQpjVDKNsKSx3qdOvt5lRTzLAITPRnB2gE3wcB2kGUXO4JkW9jAAKY1PyZUz6x1
l6mtdBk+cQtmM79rRW+WYLkyNPQsZxs3GS1Hbl31CmPXQEsl6LreicKuR3PaOup/rs8DYlm2VpCu
3YlcFEtMO0UaaUfnu33n3RnWOHp7wtFtQrqbxWYI9ebDsoiWjhqtry8V1rto200XL5QrshvRDBmx
2dBQnx6a/tlCBsfWxvkaJ5SspbtFPnbQ43bsyvp/CHF0paI60HoQLlsxEMH7OuWTKLH2ta/P8/1x
cK6GOv/pbjxv7zJHY0uNsJjv82080gggoovgrj5O9Be2HYMSzToWsL3YlQHTYijf5+c/9sbDZJdr
AIM1BTg4epbeZTsaUdlpdzhHDNGqQRlgqXSOAW4fD2xGXTYwxKaoomRR5YNHA4qXEyVnc5xNfPbT
bByKZHg0GdFumPY2YpjMTCLJcK/YVv8XBL+hRDMsadgCTVpmGE4HVqfGRMmnKnccZ6BaGgTnJ8fG
gHW+slfv2CP3Vlyv/J8UYLChNxZwdkdFJHHjchc8GxLNfJwuAyluwGUcrCmszT2LVfRvmLjfhxlK
lALpYjCN5RYMda+L4zfWAwg4+qaYXGs9p/0pRmjm+cctcQBJDDW0IE204Re8mQgGx0w7ryBKwV9g
64VTCRg3NxJATWmkKLEYIFoAm7xWE4OrWUe7jFOJUHwLBqUrk+UhutdE8qjLRzFXcUTAUYBqbguT
BjQT4i3yov0cAK66BRUi4IjWzfadn6jP/e6k0GHx2bEX8qmlU7FZEjfYYrJ+7Z2XT0I3h2r3dzPA
zP62lLJsTk2blb3NLWuybJ7KnS8MvFSG4hv9bMl4MtmbqPxQxAV+krJGecDA9T1s5skmyIJQIX54
wSCqhST0NloJYNWNYl3u1OcoL+fs7SAhFmVnf71RMXfUF3pWApCuFRlpzMy5NXVKNuQZ/OU1zyVq
6A7+cp7pUGO40Lx1QMBY9X5+r08ugn1O4Cedp/VckecBZ67zpVafrV3c0hXdw18vUprwJoXfd/rt
g0IFJfWnXaicRWhnGGoLhlTu5NQJqM7XNz5wG0IesEAd3xGAuzwmM81lYbywQ4eQrZxYoHRIW6f/
L7SP/emOQLf5xacDUVTPIOntNTzAu0ZgnpyOFFS2K9b2KElGXgwQzy/SYCPFsDVRnjxYVVoKz+u6
+YdnAHqYOh5HO3mLdmGxHUTQRB9gyk6LHOTw36AiMxQXwzrOdOXmQNjIlJZ6M/lO8YnjmoLhwweO
ZjYuse13jPInmX7f8jGYKw7pHGa2fHaXDm+UodbhFEhG1rEUqGuphKsvqTgDQ7BSfU5cqN3kceug
8fJ4KCtttIMxas+1hPDfZQ1EtIGzXSB9dOOefCulfEoUJTDHL1sCBVnRhYZ7QoNTayVI3qxudE2g
bspsNLOLLthmJ36id4untBw6i4x5UHvrbhuT3iNdadkNVIM0Kpm+bfZYcXwekWIB1NX4UrNt3SUh
GcNGlBYO+mrk/iEEVOJDWkE1KNhN9+sKv21yugy3jMEA4RWWUjM5KiYNw2GB9HFpdQZ4rk0n6VeY
GSJ/e8pWE+GWbg9Dst0SIxDLo/zw/dUpxqPhbNTQzUALx21M0tcjnwxfPi9Ow2nu3uZxyTmyk4Ae
9xuz75nmB7Cn4aq1sJcYXPSOLaPQ4089sor7kJbssY4/ULxHgqa/6vDgLPpQzut+4xY1tB5td86D
pc1NYOACOJpjlw3yJsykMnwTWDONxBWcE45j7bICXwxqRsoNJOL+AhjwQULlV88IZA8QQIRkqady
aZqeXy2Nxnq6srXidXepQr8MdxmeGzBeXMvslsybg6JYxb2NmAAhBZ5NgCQr5PQ/vuCIVxGuP0It
wX8Gc9HPHFdbx7JkV9Yxfh7yRfEN5x9k+1SvZkLoHD/GKvHSHvA4o+UsSIKeJEO/5nnw2dXf9d4n
pVZaGa8WMW3WOCx9s/HevzYYKDTXkWT7JHARVkiJLXejU8xIR1zJHI+1//kwshHAvRQxY/med8gM
KxwHqqvbZMmI/mWiyJX1P5NXNVS51Sa8EjEWwYZTkmN3hlNcRicitvImUfGxAUidrKQe2n3jDTSr
3h/LrA6FZD/YXQ7CXb0QS/H6HPBCThG+DfGVJgjWuvjJSRiX5pYajLaqIUFaBGQDdNPIkV4S2qJ2
oayf37GkXz+KvlmX45xiDaS6SpQyK0MTt1KrRslkzV/U7uCKea8JtQvfEF3R8f5mJdmnkJrSduIe
NpVQYwEj1YtbyprxthKJIt1Q/RB/MY2wiPVbDRGplGrQ5PESW7sayBMxNA7jpY3YU4UElyUXFDoE
b39vPMTIQc1/1aiZh7PCi9WbWX80VNTRX4mryWS4/exqgIxqh3+f/uXNdTzN3+7H6DHkkHSxhGr5
Kw/1bdyRq5PH+Qsmlykgu/Ue3eJUq5YbQFI81igpjHwO8Ub1QLqhoz5vx5eB/+m9SEwqkhPe1Tcr
n4ktfUP5W403UwOjBcesCYBRjUxHsqqkgefJ2cp9tsHHL/3fZLn8YHjT3YGPD0rKEtRaAgTjOOBS
xKkcc6p2Gz1e5DQrOIDVFbaT6LP9B77/00oLQaa2P3ukA3DtbO9F+g/2XT4DEG5YzZji4VenZxOJ
cs/AaUX2kOVe6FOb4ctAznBSptYXs5Evob+rviEHuGP/bUPpLWHYeYWZbsCMbMoqc0BtA+mWyJah
hdi/nhZJ4bhtmBtGb2jJGUeaxBICAEASLf/SEUCkp7gkuP7trm56+/ejXTrJkg2SMtrJn7uA9tMY
bj7hgTbYPInMpgaNdoX+2Gyk1urt06JXc/ab4+QRR9wUGIDKyaulv8Cd/oSO+Rjej4vPCzq1UK0a
Z8smpMfjJLmu/4AZYBgsKcxGMlpmcDWgBJZjKToM4/Xwy+e6SvGJIuluS78nxaMyfgwkuX9CTbBI
Oox9DSyvyqdMD3aigfKin4d0XrU64dub9VBnZHXj217aTUchXoQdNNRwoPzRTdmOameaAqK+tryG
XQ8nfIRtsC6b+kyaptLRa1Ab7b7OTL/XDepYQHNEafEw4wVKzyniNpMhDfC2s9W04dwdl8f3LfWJ
8TBxPYrBLnS4y7qI2PlSGeg2EoCimODMTkgkA6XC+k35vY17GNeYO12K9TJ+v+HeZGBsh2o47vto
vcyzE8mqHa1o4FG+PpTJLlkw8Xu98145vTNNT4JuVX8WTeFXw3Vg8BUVYx+HCbdMUv6gL/BYOn4g
aWVMAjG0f9jJVYgnWgrHs4Y7+7KyB0xzR7/VFBd2ropZYGVOCUXsWcwiSUc6a/AIYIq/4I1vUEvF
yVsEmGRJne92gmaoZeIB+8aZnT0a3B90/S/EetNpEESWX8CdIBVqZU4pR33cUJ6D0gsfxJsouG7b
OhQJqlYNABx4IWc4fa1G4aYo88ckIWyVES+k56bF1YYZtknczPDJFZ2IPT+60wGiC+j15S+Q3kff
Y5mWJCwKO0ThaB+MhFmqpoq9L+g3FHOtW5OUra5anPLf3cPaxyPzxRpP+CrC+2Vul6Yb+5AUi7CG
s6ZQPQH2ssSNWWQLeraWpUjED1Bh8NzjnFRGepIa4lUfbm3M4PWqrerY+pZbp0HVM615r3KnV5Fp
Ih0vFd7OaWaD2ZBmQUqGhofSO1hHoLuv1fFQcNWdRN1iaz53W3BL8/pQdYbOzQdpw84SiHRkNajU
qOIoDwv8XerNLud1YNbPgyoktm+gFUtgZQ+r/oq17ef+d7I61676tlolYbiImRZC7r1EKXTw6PET
EVP9UuhecEG0xjSwUUe9TuiEJ0CsMvr5NSkx0aqIcvfEGrYG6olUgjv/dcVyWEKo6puKfR3hz6Ek
YWtdjra5UydC264CcZ/7FYv+ttNprJ2U+ceH95Z0LlfzfqGe5uCA2vEghpBMGtKr72g1s7J9CfrR
3Skx61Lr2pbVSBRD+tjEvBuiD9lleQYwq2vINGQ044+nLtGUl6qUbpqgxUjSDwGo9fiDKX8wn1YU
md+39nQmkApfZNpfQO4YgpfSjmvJqlMWaydSoZjVJvE8SuxPLWyOh79CSws5AAX81fSH80FuaiyE
1GA9NZaxS+fmJQuekxNl1cGnwNc1YfbzFPesQCepYVbBxlC2yk6VRxjDSJ7kED8sEI5eLtXlfOCR
zuP1NCc0cNQvjBOusXUv2YVaBrGZ8TdB3+BW0i+YR7YbgG2tfx7ywXSpS6tpjzqliC/NMploPR/n
8Hi/e50J9Oa4rksxhEagyvs05hMJK1vodZhHhuBJAeEFkb59i1sAT3kLG9LzdtA0VN3SOlmTUyI0
FVoCGTjWQQlmyFf0lLvR1nXu5Ewj6aox71pGGTzmBO9RSrce+/jw8j+xJOwMfgHQzINcAR0lnqV9
FtaXYAcQ6pcZeSye/vVnq5v3ZMTJ6KfT3leaRAhBVBlGXIH+kjzdmTGLpbDk6b/dty6WbpZzdAb0
6gfaI4esMX7nbQvgSllAcgf86EHvuwrxCU//DGNR3ovBQl5xE/JvmlB/qbLyz+9n5Mj1DHevAhoa
WNfS87xgKpw4qNrmc+a3VxGyKTz8zI7cWwp/WldlMGsvL/LKZ8YQ6Dxp+5OB4Agpn/3wrUpKVV8x
TD8N7QYHhsmtGomPfrVQFpM6DT7djFeimFvdBjKNveKDzzx3CsWccWrubQ3S/aQHXGYGTZcTF1Dy
VVle2lo0kFo8fJ9X9+WFRbFK4VNGoA1Kq59k8ILJhMke32wNe6iFX8ATMyrx3TgCzZZrptoo8QoE
dsgKaRS/N3zZhpGWEmlJF8zrmfYD8YaHvx5rfTzn+Jt/8Zc4S8BKTobLsZKG5DYWHSDqXhyQkDSL
3RQOI1eyj0LlKZvWIcjaZVwIYibh0NMToUjFhDaPG3TiWaNm02OBIoehYu4KelgmEzXxZfLTW8ox
mKZhq8WgloWCRtZHkeySuvoJ1mpHcDN1oBw1WqWLfamFWjejaN5mjY0zqBUWzDk2mgXhkbP7XmmF
2hExaubNgHhnkKka7+C7qBrPUq++p2rKnQiznT9R6f5aaTLUPynvZpx8q8iVoeMx0VVdsGB8rYuY
aNXOmr/M+yNXot5jMWsTQx2QuiGzUoksqttqRLMa1wSKa/d0yN2hXospIIAj45sw064FPeObiGTT
s+UiPhaP/27zdAdtrEdmIPdKZhqVIf1cqfb79QqAyFOIMo0rYpNuOeK6sb94xJcRTWfYMixzn6ct
6CNRg0p1MEQIq04rENbfehmPTgay7oX+ImrwQNZCqBRsF4DM01am0E+fOtenj16CbnmHbJgoCarV
frHFsqidvmVV1U5Nd8srxeez/OOURoHNIn/sqB2XvyI0eWtEFhfxDLiQdJr9ytXntLIODoHjTNb0
qCb1bS/jsVGD399Q5dm+tXJ1eP3DK7tk3WACkz7U9E12kU2PeL9sOjw+RPhKEvq3OyBHxkDpFpFo
GNraIU+ZgR4yhb1EsVbua/AYU+2W7omd9DMBWkxSLgfOyZ1z8poTftqIWUjRaWRokpWrLbZV0tap
Fodfo6+XOtAGCU5RA7E7nXMrgV23iLiwUpjZu9wIEryCiOB8JWAqEI0gf7WyY6Zz+0ekJKlWD0e+
c7maix08I6fv6Az+VojgwTWPVN8goPkdNWHA82FeHOwOvb6yV8YcAtoOL0NQgpCFyacWjbl+QcdC
TTRuscXnfmOunpC3CzTGIHuRBU2AL9/2cq2+H14cnMIZkkIK/5NzvP2+5cL3H9YeVkhJKKvcfztt
CZO3P4v11LS1Ch8RWI6KHkEF8pOnburJPUWwzpYVarnaR4mKznpUNB625qDTdRZl2L7Fcn/KSJPS
a1vXDeeQNAe2VeTr6ekUHs/etjLqTquyJx5W55VWOpuLS6dqlk+jJihWa0tjTmozBGHaYRv8M6DK
s1q6VOBrkoTd/GjCWtnAuXejLUgJHfR3lWz+zBeilwSGo2VsIpQ/w50faq/TPxtGZjfpUG3a3IR0
YacSniKXr/uJwJ7xu1CxCZR2V8DUv5fEfqzHYnjiNGcUjmv1VjUr2YQa5PcD2r7DTJDn7HOE4sPx
QmfeRHWvxSb6UcrUpu/BG0BU2j1uBUsFQ1mbNrRvOUok7/fOdeV7vJ3TOwRmcg1LwZkiLY0QxROH
M1zpxoPXQ5XAMC788z/s3WTlhsZiHeeJKEpOU6RursRW5TNIymFuwlFEXSgs70GNYn3KL3FWV0bI
uHMHd21fRAg9iWr85kxmIUmF+E+mUlI/YSlsHZsVn96ExqVCmIocm+XHiZUhmkwKTVYPttTY2sUR
1jj/0YWkf0JkjZvPtoz3XDg1vCOkxn4S4H71JzHm/wZVJYmr31r5uMKaiYN3o88F9F4klhWJdXjy
N/N4TwJI+V6sqWQmxLLfjbjjPLkErjIC0w+1NcUvO7vqUNkHhwkq2pYPbOpyTT3zeg/5jRoEg/Ad
eastWhrRGFjYikIxtSRhzPP1exrkoS6MBVP1XQ1TAh0E3S0kxoPqmLuzR2lcKObo+J9/Sbo228rE
qbHtaalYhJ24JvvLAasoD/S/lczCXFYAU2A1zwt1tokrKWs3m4zuC1+cYpP9mbsU7rJYflqSxdXt
e5NaJqI7zZhzEDTY7PacVE8rzpnm93i8scj6DRdViWzhN1QIDvIlJtZzD/uiOJIkYVfTtEdsirWX
dmBpn+tFYQPWury+KbLdNPjyoS5X/eGb9yMaPHRdmnacuFsyjhEe+WOiLn1M4YR5MUv8T2ftKwEW
FMDqDcP1dg7sR3/9tUF1tNa4g8XeP8jTBlXqg5bBjq0SF3aCt22PMT3YvTFTpV8jAPgf6yEdhRDr
OViSwrT2u0OAs4oqL+BJj3c1nprNf7HEW9+XwlehT3x1GSW02vPSeGxUUn/eHCAOTbk3YvYy3jUo
3pHPpqJdZovlOuoVxeCVvarCEPc1FPR+fBbVuFwI/s2ZeOCma0dchaayA3AQWvpwRRWUtsg0txVG
5f+L2q2v9E2l3PhP9L/TMBk3Sxhv1pJ4anWanD4GpEuerZpxDRHnzZZrVtiiP+0sgp90pNIeL6uw
rgjaZEGO3O0jm9rDS7unl7El/z3i6JSKATvuUNZx4brL+oP/Wl4e0gaW7g01c+X1FXxwAAw6Tcpv
fYxe2RGRyF7rWE/56vIwmfktKJLycbB4UV4q67YgIteVbTp2PHRrQUMwfdac2reHvalB2icC4op3
J4w46sCUpxijSEATNklzjMwDO+fWjeWcVokS4D1VFEHLElozlADPO0q5HLIQPOoeTzKfb6DnFUFs
eksnANfdhQ/dlWO8y4aMy718MY34je1of9rw26CNj6W2Sd1htZgFcp0zQQGGHbKTigpIeAeevarl
hx1dspEerIKYQnkDBQKJp6O3wGMbfAzyrOKc0/YXY10O5S8KY4GiBkHBvZrz6XQG4z3B03r1nY/B
ZrXXtIdPpauZPxLjAetbO1Z5dPunA0yiprMqv6M2Yh5hkOQQuPzHrNo/oT+EJFlu5ei8yg6K+dZl
q3D9rmE+x+tHghh1uf7LDNCpYlKpLe/EXi8NoFb9OJ6jlGvA8FO9TjjzQHSBQkoNTktUZK5dOvfE
p6aZK5SCSYKwzC8XMwS6cUa/erQ1wbr0W1OcvANXNaNcmZrxVgfh5dq1BdY3ewhZNYmCC8gFzKyo
E5Y8M69ei6gQvp20/6FZuHA7Gc7gQvTrY1kr6423Stfc+730B+ipw2VC3qO+JnR+ffME5mN0p20d
WpYnLFSDGSiUPMeGOii+lnsGdTI650f2OlMCYHRSIXhHEDfHw4uWtNM5xDHnDhgC8yqyBsYyvnHS
CC+s0EmmGDFLjfgdPKudOIYrqNY3uxYfH7poYSVhuiuQ7E7oueUaD2/I+9LjfBo2JLt1TeCA59ac
Jf7rv5rAY0OWLfk3EdNf9Q3ivqc8U8z/i3dvr905/vV6GRIhcsisRNnw1W1xVQnt1yEgqPUmuya7
sGS4x6N9uX1ZtxDHmsNhq/KVAHbtxMGAWkcopy3wjEHqRx+zvnBhGBE7dsC6ptc0ZmH+KV8OVLbA
8MIZkRzL0bftt6cx5B76yUvWJG5cDqoRt5kqTfKhGFGBHITOi+1l9ZispGBWS15RM3pYa+FLaQ0o
Yk2r9nq3mMVtDHqGWJ8dp4H6zGOOkaoviOPa1yVVc981uajcofJ0Gc62QqoDLyh/ymvn1+a2cp2I
OoLdFNazhbVNqCXAXSpmjhdd36n+OgHCLnZFg6DQWWpUV2gTdS6fWjNNOpJy0Gc3+sFCuLimtweU
AHlCz0f3JwW5eKVT3IuvJnGR2+1VdWWEhBPb0SlTkkSHWglO8LziaA5fJllwwwbSnxCJTuvk7RaG
P9qmEtMuOy4pLlZYcYTWywHbIa/MjEa3ED4WR6+7s+37UhaxgcC8Jk/3SW6Q/OZdbO4fDU7sBLJ5
YaeEtmGfbqBoBFfvd8YTylmrWVmxqEbDqmtaGx5W6sDIyqJJgPUhT8mQBvGQhnchA6O5NT0ujNUh
h8iYb86yKF6+3+x6MXHv2aGIsbckk5XgXNGkPAjcNYruNaxnWANuJ/A2PqCHCbr4Svusxe7evUIV
ehcvWrz4gtKGE37fwOd4nRvug2KutGTIHCuH0yE3xFJ1ncfUeDelHSTunyn1YBcDOxLiVyu7CZai
ks+a6DB+5X4iqaeG8UO8zLW2YR2isughdVolc2HM9HBspsA2Jlx8KobWq70OT1HKgPbhhHthvWzJ
1LBUws5pGnau7rR36/cgVSsuNPeLm44SYqKGwTcgBbNQS8qSmcxQGbrXtzlrGj1iQbSCBa0bzz0W
/ArrINLOXZBpIzHzK7Uut3dbgcvQh+up2tbfGF2TrZllalCn3SBqEB3+RVuudQGwsjSAkVN1xzm2
RUkD/JT2MyIYMRQhot/wvhNv2ZBJFiiuDm3fP48pdEvyiQ+Jn/uQzt29IgdoaQYX3Ea3b/lf5znd
FWEvZmfnRpD6oYqysY6okyGaACr0oZydqLUcLEAo/WolmYlTCvHtgMIpwhQ/yDpGqJYx4T35o+8c
1PKgft+vbKbgZU1EDxLkqcN/cxTPCNdhHiC+c7iSraQB7mReJNfeNY1PbzuwR/RY/jezLS04sKLK
C4XEdnB1M2LJvQkRtEu3d7hJQINdzRe7wChoNzWGElSau8ZybIkFAciWKQpgKi4C4nkMoTyMONvU
vxvEs7Gcv5dS7TPbJ1wyQyPCig9oP5osgy7wYIdGORTuyPdpQ38mgwXlD4GzL0L5hVbB1UOnbW/K
5pWuo/4bbvT8B41JH3GBp5/PqezYN8kP8CegP4qt3eJarrs4UXXVQGYQjQe8JCcFjRL7FmCJNF8h
uGC5PwJGLWagBbhLE8EUo4II2LsYS6CQUB+vPlUAstyWxkz+erPb+KImUhdtxuSuVObhMeku2p3o
N97i19NTKWh68npdEiiZzQYeyrJPiiUfApumM1hE3mSmnU4gPHspkYhNhb7ZxAk+t5H7ZHfh6wUr
/193LKYfsWikPtAgkGAMqdg32HIXR4Ijf4h9eT2VKtAFU/5JkbEwfdPCBrkVH592HDxvK5O5zUUb
R8iqqVL4RMehjP+XXTbB9NawZSiu3UA6Dn9LwpYquNx9emTkEhROjQEqYxX3SI8TdiGJd3KRehlU
vWx7X2hhZUqgcPXipY2vPD6CEAL34LBN7RWDG9zFuYL5bcxnYoY7DurWGwW+Uu04qDZWHKuDtKer
1fEPuf3qmR9eCWfRtL3MeWbqSEHmxzOct645OTDxgFB0SJsHV1ZHxobHJkJhC9xkKLZNbSQSAxpg
+ypIIs/1/29oksNaTgDc0grk5lcloY3ZqHqsEJuvg168dBFXAlREHDB04giMzTxbTfNcBmA+iix6
1u1535X7cXu8WgVi2AKpg6+C6a+YtbkV0xu42ViXHVg641gQO5J1p8x4WLBdFsfkIcInbJ7a0/bZ
Py5bf6AoHg5QMolBbPo8K2fGEI03i5nFkBBoP05CrBCm3r3Ti4oBaWWog5+Zb/mEC1Ii9bgCvy9u
ojeMwHDn8xrN5cFK1dOqo3YBlXGMjGjk6QvQe901aIlS/geHLU1lffsyKl/Oef8apj12zvQKqlow
F39RGYkPUlzOTtW/i4qdGy6ESAXFPLTyDlNGljAGsKKas1iF3df0XIL2G/3hIzRFFaT4Z5N47HAs
EGiJtOhQ6bFPpOj3rHD+fceGFsjs0LYkJ/R4SBST78Gjv7tXjC/QQ0LGs3bzwTUyYpu1E/SC65F1
fUbSSmvyWqs2CwTKxVH8jzhWHK3s3v6p6eKrM0TsbNlScPJPRMPw+JyInpTrCu/ewSLJC6TVox7F
zBxIs2mhT6067Ia+1yeGC7RuWULH1Ybs4L64pDzzU+T2LUoi8OXHdaugPgSDOKP4/f2HKLC//IlM
3PndMtN3CIL70KWy0Htz8+WeZlszOuruCy8QQGwPCvjoR4rTdvQ+XJvivHrqucooWnB3y4iag13O
OsswdyF1owEcjs1N8/3iuhqeR7PVBPLUHuskIjAC7gyeQWJvrvRrgkxdviWqOx0MfP+0ouqttPC3
eItvLqGu900Ssz4R6eY7Z0kDgiZn3LTcNKdpPkHxLZVvTxNkv89iu5CeOb5/CoDXdukx+80Q31ax
E8uA3TTzYgpncGt/tkecvGWckBPjuAY+lBTXvn6WpDmBxRKZ1XBKqw3ASgZk+UUeRKz17517v4e5
Jogni0OziBxZGGOYwswlwSp412PAejvnaNEtVKglDKRkqhkzxnMNtQeoahDvLAKdwOB5rJ2evolB
fDKhOn533Do3RnOmLDWUBIUdYyt4lT/bIsLpKwwhUirnWTfYSslxuwvtmif22fiSIdmoT/W1cNI5
CEF3hABT2fW+Vfa+58FzCxQYUkx2ELHS5NWhQs10Ft5tnuf8Q4kSqRzBrlEas7i7j2g7fuaZPR8B
VvzjrmToUsfzEvSzMfHvtnQ2VIGmGDb3Hurf0D9gUYMIhuFMoW2s3OPIc85+hbw9hdNVT+SLpGy5
SI7zpYP9hErZt2/5faJa7xW8gaafnQRaoxKpFMwtVxfkn2vXd/rRtaB6Vw6mBoJMqjkr3vX+Sy5W
kwC2390bdPF3MVDnp+5p1FbiLEibBO2Hdyey03M3xlD1s78c1CG7yIVv/QhEuVdpJ2+6r0MOL7zG
S+35K+IzeVHS91Y5qHoS41lNqex/Pvp3qqA32XjKRBBNcdcJ5pyWbGeh5G+5ohbfV/AXVY5YiVA4
3H7NK6me4gGSGeZaSjLMYV0k+KFcFiHcf/yZ03QjG6l8OZ6quU/Ffh41MC5kD6KOE2x0BJWu/kO7
AcAYKGrk2ET7KPY89kIzyMtIoguuygEycf1L/9bRBXXP0Fh6x5IV9/twc24Y81IhvJAo46dWVTrV
CYPuEn0c6VeRPIGM/YwSy4KDaYTnb+/xFTY95IxkAunip8XJkmjjeKedRpYa422rUxcO/zopRogF
CYFqC4Kr4GWDTuy+O5xFMf58mj2iiFyDhUqTFJV23wWZ1WU9reUzfORMSBrnqO46xxJb9sTSpii7
CuRqxzH0jvawG+o8TNeCv9fSrgatUgDLMV3u09Rr97RruJorchkV5XSvKSm9akZPnQh9jRE/obSG
k9Llog31rIVP07NW7UYZhPcXAI8bCz6GyrQGe/olM+mNR8+TrGXY08FviOJhJ0zs4NOhrxh7REVv
E8T2wlxQtLqgoLN+1mwbquHNq7OnWNyimt+Xowtahth604AFqZQM4p2B9v0HqmH8n/HnzFMTqPyU
RSCXblANuiz4Ika+qbFfEpUA5I3WlgyPW+1hqdt/2aNwg7l7CPdEN+FYAR6SuvT93rX5fBt2V7R2
QJrJJUrY5bh99YYesNVwV6ky1OoLaoQZGKcP9HzML0BFyYpCMg/Pla3z/CjAOiG9+Rx4OCavq7g/
RcOd9XGnRtRUc0JK5t/CGeUWk4+m32UvuGpKFwMIMO/ecoK8+jm/zIpxsC0e0rcCwCClOdjeuuwd
TlYTkes1fm5a9WIqeoQIu9lVMibtZXbYVRE/aYjIRvBh6pgxDYuJHfGYHMeU/kcx0KKmqFMD3zXE
6iCncmZi1ypjPEvrg2aJrgFz0Eg8y0HMPQkgRmXzHKC0MBNDXFBlFRPAY8XZXf1mn7kEAaMISCZ+
eUx4USr5vJiw+VGJwIcVDKEJF131bilLcYWwJvx+TU2S4yQF3u608osGrqH5I5PQYWisHbz/LZNM
63GsmFq4NIaJvSbO5DKjqb7HPOui0e2VSrd6RSe4Z1p8leTWFq9CrFj3D+1e/Y6JFz/UxKhdJGXg
OImOx7hLB3t27XLmGF0DZnKi6uXtyd5X21LXVJpADz83/7JWzVc3Cqa9LqBxQrbxArLyqlMjycFT
fNtpIdAPper/TW87XZftD2Z5mGiHFuuYaWvwmqqvQt4ruSxq6E9zye/v2IFyQWy51ts9FqV/PImi
zmi2zdRzvM+bAaLPlfwJnswMeETinEuaENOZcM9is4cGOjOVy0REVEa31bii7BDfh/CqRPOxvz9z
kovQZ7SdYYvE6kaqHRisC3uO7XI+8Ovl9NfN9GhvaYU+76fjTxms69moBoan+UaRILqHGxC/s4N1
WA+jiKeP+l93I+Ii5KhUJwQFowomXL2kbtvLJY6A4du9ef3jdRccgZAiTL2wwZIpUINaF3V43FPG
vZLTCV3W0FGsQH90lqVZPBfR+U6bI5vkB4P8+ecGqgrgVplQ4V67RCMobBkT5E3jqc1V3mzbmUOj
AvJ7i0xlkGLj49rTfSO+6ieIFD9v45s7K5jDQjCOACZ1hVESzRbIWWOZHin5k0g//sorz2ilmzRG
6jzVnyA2iVnmz0YNarRx5n2RelCWLEChJnhY04ntl6icYnjnyWexbMl/j2Pw/CM+jJgbJ5b572Nd
Iz1aT3qTRhh3iUwTh+bLk9r/X08OrvKsMQC5WvHhWh3tcdYosUPVxFPtYbe2HnzStxYg82ZmGivj
N8TIS2C5y44EIOkvCedqwgPimXepFgpIPxDIXCgL/wioYPtLkmGD4cWX5Fk1jV8sTcI6FGcCTkHc
7Od6VL5Wcoaome8jUnGWfondbCErqP4k4HywMpN5p3MRzH2AHdXTY1JQPHVlXgapbv51O42JwjiI
sos/nWWA18PA2XwTYa3w+gXo/uH8PIoYyRbp3cxOjUZY0hjG4/DQjPMl0wSLqwaJW26cOyLTu29y
7CncHE8gLMi3ReKM9JP57td84UI/Wi8PESfO1lxqztQ1D9Lpzv2uAz3NmkGfrG4zm0yB9WC1WPzs
CqAiQfZI68g6Eqk5MnY4UqJM1YnRj4R8l4QfZ/r/l+xy/ehRL0pbsB7LuqEzfA4+2nWK2wWcvKMI
egBkICjQoAhPhoWCFVoy/1SzZhKqS1LbUJCvIzwnykCfoep6OOMIDsefscfPlobwtQdKdFx6r2Q6
vEhW7efeGbnahG7O11xa9nxXCTK5e+NhFzQJSQ51R4Bl9IfsORE1/Fa6VY53/CXwbIxifMXHykyL
tGzrgGm1uR5OQMF4TzFNQqS5JwOopL4cACpZcD6eVwxzn4YoIMR/mGEysu/R+CBCAdc4LEx8g1gd
uyNtGlJzL6F9ojsgf875Q6tJSPuWmLuqCOEBncHiCG5JDKaYSVljoeLjYDMqI41EhwVUEOpTdVhJ
F6tEErMd51SsO+J0D0oifxoRnjM21Hy2yNr99xIxKVhO6qcdR2v6UPiUNmjKVtwAey8Z7t6lRgxW
j5O3yPuRF4uhiTBMLAU4e8v/TmNiM2/tM90/T6HB7vblj4xAWtCIpOwxtKvV2WxZlgsUq6s9G53N
TGQdQNjBJCapPqcK60MR+E6Jilb2dSRZibKZO7hxk9KehSTFnDEs2Yk1LuuoYWhllxWuul5dupdP
T1w1n/WiBbUta0E148G4csnLYHfn4lhkB2w5Bq8x5/NZUy9UBci/QZPmpg9TMZup06nQp9fABZtX
KyE7ZLjnOGuVCps45GyISnSHcC1PAmpWc0MbKO7CeRGkaRgIiXTb9nTrrUiFLMN5qbyCo0h+HMxp
tlfsJmJEAKYGLC5CmQORZt1itI7qgOaiazUh3y+KTGhNnPNcKARUa6QknNiIvqCnxVfR5InkxuDB
bdvNLmZYAr+ZaqSGOIbhjqLgghH+ILBc3Vk3/Q7vod0NFnxLQNVTPJbJC7ZiS8ngmGS8ixA/WkPf
r3zvutMLcy3mt9qVcopnEUxVM5mH85HlR2xF+2XQigS0pTomPIJC6tWDrlGbpTHCMIoxLaiTt3/G
H9UP83/dqL1+jUEVWKmJRb9CZp0NOCrauW1jOKYHKLc82Iqym21hydI7xfVS2IRDgQaF3vfQSC6y
fvw3hkae8TAo9awy5EtXzv9FTvReHicGYQH7fvs/5XQJtVClWqStC7qOoFT1PdQegZwzFU04jz7V
EaqSpTXoXaMGRAkvZcrkXLxwa1MQa1KyBeJzGgg1bzpXVMqyjAy4KvI5f77RFj031Lg71btwJwaz
ZbgyUU0GHmm+v+wcrozcPLlnFYBxhSptG6uykJyu5wMqdGFd0SDiv1QJuDia7aTpdJ+cVdOIBHd9
Nl3ESylgo8pAyDXqGzHTBDRcwf+fghjxKFJ246E8NoEJF8/EJQO559EY1kbIcAqHiSRnUi0hoB5W
1O+DGdf/py5pp9vLhmwUrL3cdD6FQZ6pecwbbbLJAfZPVtHbJe0Th6UaY/J5sSvW2jOTLoCH70za
K8HfQ/SvYxzVKqt2KHR1lYEssWbrBcl2bhDYdkcTHjH6ZnpAM57xoKyv09RapFMQFLD8s4gLc9hp
VKiFMv5xw4LuCt5en4NWlOQyi1KPdgWxmQUUrYdPVCxd4Dn5rEpSN/0vn1/b8p/5wIS9LFhBM5v7
tmF2hFz8J3RDszU5PNWWfRbhIAMEDFCFz/WehByF8QwOj68JywJbqkevRM92QZGXov0V8f5SvrZq
1sXta4M0R579qGw4mPwf60emZvEgdUp7NQ94BkBmcRZO2AfutIfCG12YSc98JzaIdMldLpKW4E3i
cPngRZt0Y9EaR4LWRpb1lFcO1/8s4rANHbboQamSmfk2rlryqsTIEIGkfBrzJyvfzrwqp4R57lL5
mW8w4C/38Sd3hkYtKCFGiNK/ddtT45O98Md2AbW4+0vcgAkWgK+EMcaaDOFOaFT29WJm7DB9gtHZ
u1pYE5kWY7UgfbQzROX7tQqEDj80c9yEqBfzEdnLgUNenVrlP6gkgcOabLfNr2UfWBITlCAAlU8+
Ue7TRAemTACGH2OdxhakvV2n0oreQ/mBjON8re+yM8WLf5JVrqWmm2Wi+VWqweZzpC2kBS5gsuRb
BUhvv+gm6593Q+y2UcI/mrdRVFqnF1uLrhhjdk18+7V3k6l/Zjvl/xekAWWdeqMZ7E2r3TF+6V4E
1V6P4nicIKpGdkC1HgDMtdsCSP4d9YVOSzXJnTP6+jPFLyuORoXI2g/XDM6ulySgHgkAh+Ryzrod
J8/cnkZv8vBvOiNhQ73LxtNizTOZD2p05UG9W3tFwG9m0dnKXIfB/wriafJsNt35uJYBTqD4yCJq
Yjy7fKxHh+bqD6aE6wT42Qx7P3MxAd/YqTUP4C1FMXqd/F2DZQdttZsdWjY1q2g9pq79Rk+nC+Co
tyUuzc4aMKHQZBmHVZH/OgAYp36Jm2z1UTbJQmYBklE0m0iTNdiZ+J8xln32QpHEn9GSYOrdb5y1
cepLxuoRCdZf8ai4Ox1ZZp1x38bXilPcOGS8AUnptAY2o0SKh0nX0GiFddnot53p9pIguXcaxtfh
ElI9S8jH7zKX2CRAOa10ppV6VyJHhWJkPbmKUjT+cYjz7Oq1ZbMk3SHGaLyICL4uP67g6f+J5Fme
GNTyNGbQIcXYjn2CgPI64mprCLOUEkqbdJnlGLeylFpRrtHxSChgfoW9bF1UhVUHgJuIqYppqAtE
CbEutN/IA1hgFSWwO/CTMT4NOWoJo8VzdytrGLpn/mJ/1Fove1Vz4Y9pBUq3wqgf6HhMs4V7gq2v
/8Eu3OMf/zyqhyTCp1XTB/Qjq+iK/oVtdvAPnOr+VN+6x2d04u+JlKfiD2frMy6duibXuUd4YjKy
yxxOppqTRezQUtRlZeHiKDR+r+R2gZ2+FPq3FMdgxk8AEsWmO+bCANlry+8bMVjXewahnwZBylr3
eNLEkDZAn7Fj8+UgPW7TFk9eInRQXOWeyf4mzuQa8rZD7WVowuIowaZKrJKk3Z62O/sQDf0wLKVQ
nTHJhU5aM+V5dOY+QA4YDV8EQn+1ESfyw3md8g8FzNo3mOKbWYto9j8hzCOOXEbEP3yLLgPCzLMb
19SibsfA0lYiyzCzHeB1EpDNomWgikzcf3pA/U45T52kDNmBRoH6GXciHDq5iVykgHNzHNSNq0qf
IqLyULm4/aMmu1cwCiLL+gt7xKNFYewQz2DDDVqEtx3tmYs7Nv7kLud9k+sPefKIdknchNpNKJTm
Z1C0egX988dIiOKszP/QUSKe7vuHMPo+vjFRYUSvWbmzwRpzOKqgKVTRN2eQ5++/fm2JFXKXcgeq
rH7a3dk1v1c4ROhiChAx+81QE641+CKPa0ohxJO3gbuqMMeY40tY7PGnT3O12v7ECJZ6+SrEfQjT
74lWJo9btYN6wkRDuuD41hYyDQspEu7rdQZB7gdWffaw2g7hVf4mbx6g7i0ZDYxMyeryVDj3UMIF
txUsWSR+J4uYCzaXtGJDyMdwX83oanXuc1f9gvyNq+leEXJxMVspxfOsND+KX/ZMPm3/inVDxe1X
E+kasDeHtS78pCnUZeP7kwIy7B9GFUO3oZ+2N/wMwqRfOEfQNaKJTotKVIyNZAOmsMH0uqbAMeiB
/nisNH6bJTC/BMj0PZC8iBf3SoRVIAM+IiT7DK2nT2UdBdWSmaCsjuqN6nAMCOMvXM54nJD2Ze1F
vB3qmh1qT0XqYkEZ+sZmYlCrDNmM38N3U+Ytuuvo7CQrZB6gf70rDpIf47wHNA61AmwVtVe6ZT5P
GiryoIkQHOwL1xn9ErDLGG/Ui6o0WMPdtlwH6dDzaTTXv3V9M2/oQTgJUsY04QPdn5uEolJU4Jfy
m+g7ZVuzFR95AcwkPLSSZ9uqQ+pj7zEQLAZ7mVSfyRcgU9mHW5jviYGf50UFLFANQNMxVsQVdLmc
KUTiG11U/kATE6J70W27Lw1lLN6/5g3/sWO4aFCOMYnOEKiNKsMTb48MLSbYJlsGNdAGM4HluQf9
K572sx+81MDvg4EAPdSMPNzHha5RIg1jaSZCVskexeESZehCixmvaFPF9VM9treA0gRsmzTcMNw2
oF4AQ6STaJbf+1DmRECLWTe4c7/4honKMb58ZBMEzCga2b/hS3Br+0A/UM856AR7IIOMeA4ztZG0
ntDVI3xORI/qIc8i3j7GZJo8qGYR61pc4WOKxWlPc5bp1fxICr6yMcCejaiuuCSaONYgiEZ1arN2
hA4lDoIHSlEkTYQSz4SjGSqmXij2roZ8pkHRZedtFOD+GtBRFBIC3YVF/W43Jw5e/rS6jHrgCKmY
JNxClDFd+AWi+zm9V+Yt0pvblTWy28wQgRxlOCWjT7Zx2dTxoHXH8sWcMP9WdN+BE5D/JW98DHSm
pT2JxvxqhKZL9WWQcfsknDT8LfL0ONXFX2t6wXhkQage3ebEqxRjyOUcP/fYDcgk2TJfUWGpn741
Z1+pNDY0XLF/rZILFpFzkehKWz2I4JCAYmBfz35VK+lXuWDyJcSEbHbf+NGz4mcaHzRqLQZ/58Wn
5RHUvhIYCwt98q545pO/O80wYihUPxsZEI/Es1U2OefHmCjcgZvyPR/+kk0zaU7BgbpLGebfJVUh
7m38HtZGfpqP0tGrkt5GVCsxibz6x2f/VpLNql5Pzo9YxVHgmJWjz8TseR+6SOpcomPtI8oA+UqL
8WkexkAjYAuJ0rfr7wvzeUv2HquwOKVg/R1HMi3qah+qsErnT89Oa3wuKcq+Vr4sDfVbyAf2KkMB
NPhiAF3YFtgVMJVqRwbT4MNEZQYSUhY5QgkFTfbd3DHIDMSS5SuZxzNJ8L9My4wSF/sVH14qoTzs
txkSFg4pTiWgnxK9AEx3b/qL2Ck0DaTzRmN5tJJf4FUnxe+smkt0pYMvCV7RBNbOPuBijlYElvqd
VQ+np8MKVxUM286JTyrcpKUudctDQ5ZZX3trp1y3/dSGmwYTObrpKcCXj3yjUdtgXzsVGtxhupf8
Gi8Is0+GhPtaH5U5SZXaqfL3ejtHuIyv6ej8J1H7oL1435d8aWDQ+zaZtVbEcaPEZDkqRp9sp6uk
EVISst5BDYAFwXpKt/1AHVSyA7GxkJT5b+bDJuqTiasJygCQctFfx+sesbUTgXO9W52OnwK1mksj
hGW7sHv05IGlGtUg/kod7d+/XVHrNijTGOh495NGjtWMBCsAXiPx8pT2BMIgj6CyJ3FJHAcdyCiK
OefFVerEmjJxRRtkN7p3cujf316/qq/DgEgLpn8grNsNOQ4590ct56q5J7/2mQOvqMRHgKjTFG9t
20RK51hlCVzlPU48u9OfjH+bFHMe469Ix8ngAuAvO6fWdW3c9Nb42NMZ6oaUIEki3qiVvymwQBSk
ZKOgqIwo5fRM9DeQST/QCD8aHWIsCn2zH2yDooMhUjS8UfLEAecZvtV/ZjkkRqQGTrTRNZ4bSScz
+DgccWh+n6AklBHygEpXu2h63heVl4w6C/fesdrKryW+9HlB7tkAERQoCO46bRlVApKo++DxUtW+
3gSyqB5vOgKK2zli+a63Smz28iKoOOjM848yb97vkxxBfeKhUpqr+WPC9mH9+5oLLW8CmBcfEvTg
PbmOorubBuFhfLknvO4+ahf9ouHtQaW3h8UEoZCpeFfud55pECMfPf0OF/eJJoi0FemhIU18U3O9
G6S1Lekpo+zb0F05TW+7s9f7sX/Z2X2HHlz9Awn6ahqSDFxZCPt80quQ1R93AZWl11XZ9TYdUEFk
y2WqYt0Kk0f9a9RKHBEC3brqj0fI4z6ULqainf3+J7aEr2OeTpQ9Z6kvkonzaUkh0He2fCe3JDAk
Sf+m5mjzskk/xR54WaVqVM+JIAQkFimCzGUrfgmJhukX5uoja4bt1BgA61XDVW+4su1Ryem3mYTX
83xVq/nvGYppefanAHHYMcq//Otlw6SWRw9mQjIXVnKd3G7Aq7uncLlJheJz/5jq3APNkMkhoIk2
6kWEkXSVUzsOlyF/HtX8oNwPkIGy4e8SxSH0dtHJV7Ew/JJzMQXPmKmBOT9dtSVgGzu3hl/A8ACY
+qWMU84keOC4SGZIjMr+XBopdoi0NvCvQ59CEfnNvnTvADbvWdFjXWB+Lt2AZ9edTVroE+VNiSX0
2H+ulMvx8krLJtazXx4PrbI3PJWJ+jckGjHKeEmBPOcUgh/w/YfJupx4o8o1Nw//6m/t+pFnZSup
Qp/kxbSoa6NHldtmk4ZLSt/4g1L5ERbgRgaTW3tR+YFQ4PMqGhlLAISBQzlbP2Y+3+IYZv9UXAhh
tjBrngYh1zE67T+/T9fCf56tTPfIpY0kFWpyntndG5jysG6kj8jeg8roplYIVTOOFP9dzoQTkRHN
Golisf2+ers2I78rLO9PmstwMyQ9Y1wHikr+wdX00Po2dn37idwljCPFkauRNtAq9eqxUV6K62FV
RVLz6NOVEhfIsJuohybRITZheGkPuDIJMKMUWdk7ql3oGDJ7veIB/NoGwOrPiEFvaVvXENU2K6Kl
ZFuzK8MbpBZYEzAvAqIh8Z5Nn8Qab9jPObI5kwpIMnFICSjJsHdh37F6DAk6+HFgKUEakZvJ7yWl
WfRZZXdT8wZW6hmkjQHEbrmqMkvlO/Daptt+/7vMaMDWSz4Kn2/BQftiohhltdzu8yryLeeSa6G6
5Xjq93agBo9WG7UzR8zJokcJIt+l/zA9KlftORni6vUoeQu7tf4jCU6rfT6hmcqHaQJrbSDEnPQq
varcRAIGR1HNNX6Xp1Ajtc8ovirna2K45+lRbBTeimtKUKmzq/RCJwkqER1yHaEEPvG93GbDONc9
uqSbhKpRPuzVLlEaHQYpIYY04eyAcTYje0i0wXX9VfL114hDbh25bsJA+snt8ZZ4eR+b2m9MYE98
A+Hbc+YyTcCP0FMkiI/ypwdh8mPhPYOPAiHMkfpf4gE3M2je+d42/OJLlqVZmnfbOKjsO4MWmrw6
E4AHG4TKka1vLV8nTLmocH+K+vEnC+z+RMe+Ol2ESo+pMjT/tnWbKhD0W+Y21qh7VNN5tEnqjhw9
mjUFDBg1GeaRWTtrFsxH7pB1e1/6QKWzxQ3anTLrY33XBpqed83KaMSAKd1Rsb2C5V5ZL2dF1N/Z
VNUJz7JenozVnq1Gt2LV5e/vITrsolz72OhMvN28Ja8JBAnpaqPSSNDLX1A53TgbMCHCP5ZzET3B
sEqRNo3oSuVYXMw5OUOmiR16jV2GBW2VXEAup0ZuMTlk/+M/G6Ck8vUQFWoexdY5TCmTgrJ7SFgI
hEsKvc1SnlFyvbS3lVsIOwD3kz2l1Paytjo5sW34tcd4ZvV6gB5pMQvFjy1HR8BjYIpDT/BnPDtW
8yf4M7RBiO6/MFw4vbo4+i3baOVquaAhtPE/9d12nsjWLTwZbh8dG5CSLRqtxas8VRlH4qwBXRoY
OOa4DobXD+jJIklzTBAg4RBqUptwujKi1wP5w1s8XTipFTYy5A/6yuLMzIeXEXGah70BONmdJ9yM
8uBQYvA/OO3oRx6coeYCzCtVLPWeAOnkzbpVne6/1tPCE+drTjxfcXwad5kprL7PIDgt7iYzSPYt
cA5fBdoWau8nHUzjQBoGNfxn9L8S4jmk/FdWoVxSJFmbz8QfTWxylqX5926Klb0bh+vpxgC3dtRN
EvwWz2DVg2uCA/7EFrhj7fgFExMhTtKdn02WufvIneflFv8tGdTKwC/uChkIK7H4Rc8EfrApwNUe
+6nherdMwwQ/jC5/8BXwepq3cBOrYZCyqEZGCQR3V++PjN1GcVRhTo6YUShPp0Y8KaY4rzoNovmi
Si7Ajmbv+HgBlJaQwj2Qd3BHGVTPhzoMgfWeICR74pYwD3nPKUvRwpVVWTXDPYpMEU7aHVPQaZnR
Xi6S5BkpyVfAmfBLxHHnM8vdimy0Biwf83lsqrdMTJPNfE8+La+BjzoPgRtkRCtysx23jvW/n+Kn
iOWf3CdZ+Y9gR3ONizbMK0Fke1dLhNvK4DP1eqJtg3q4ejQ6yvg8ePA+AQiEKVtUg1ihTlxDe8Yd
Zja0R4SzNEPD7akgrITH6uDWYyArQ/jLuqrPPIpaqRiqN5Aahd2Kwh6q15mlTm5v1J0NmXOqDS5o
b1bi2or8cyMrUOco47K0Tc1+UOfLwPVt0dIAwL0PdB2WjSsDLfRPjn5hVqnFlJ4a1uk7NskP7Cv0
uyWlt/pnpdUtvrl6y125GBGEVCmUAgewFWbCQapp+SrodFDA4tNeL3AQTJjj52DW8bi6OfBn6zwr
IhLGx0ri66cWmypYnkbJ5niZysDUmoU83iNUVgmB0Z/ZqVIBgcVj3zEZ3P335Xowb7qFNmtx4PXT
vXgLYIUNc7qxdWQIoaqTZNJnGGCsBjQE+kiAMHclzgLQialhiqKcCfzewB0JoYTG4dAUQDrGqf8S
KyWoY6kbr+t6CouW64W2rFpkyMo/k4GxVBOyswBnfHJAytirwq3uEuRpB8gl5jYb/1y89IKA518Q
jfjNq9trznrugF2cTpkNVrmIEw9S2QYdAopx/Y2s6kOil2r6XEw7cblZ7gwsq8eX6vpYS/Cr08EV
4H1WRW9rk8Q8Kci9zyevkIQOr1Uy0Kl9YUhwBPgCG1mPpzSznkVTtL4NuLjtDiDOFFymV8twbM5M
XoIgmVV6ERD/h8TzWQOE0nvpO9tm+8ftYngMWMh7ryhlu620fKmB5Bp91vhpoLebZIUw05U/jMjL
P2V98ZC6SUxgO4jParhACpA6mGwyO3dwTuZJDNS4nX5vvo9yOt2h4/NyO+QOLxd2Wz9Mbin3Zb0p
6YobIXDcz2zOXld5Gi3+3q4MzFUFBRdtcoK55v5rHKbqj/Xydt9NPVlFz+DveRgGU7QtQzkU0lvU
rrkIZX155LIMRAd5gL8K3HcNcsUoVHa9xmUokyq0d3xjIrbH+ws4Pd4qFfalidHau9DJgoHTG4pC
/kycFyJIJsP0RCLnUj35xn34Hu56kseTbWw2t7mZHl94psIPdA14ttxydHb9d5vOtVAqFOt5vlb/
jfNZO5ZfcK4Ath5VP751ANl6Jh7uDAdbJaVE6N4LcCjx1QCKvT0g4aiKZOnNUia1WF7eCZBvIS4L
NpdeZ3x1fEn29qj42HaKWw5AevoqdA77c8bKEyjfzS5GqRNuVZ5W8Sn/sqNa57Iicifu9AZGv6/p
piLRn0LN+PN4z0aL3C9rVDMN98jGWhkTPkZnC79jPXtSl5nO4Disomb3UJ749OPRUMWATbCWCoCM
rmG5ohSdn/JhCPeKE0qjkANOfE2jlN6FOFkrjI6SvyeT8S1NdY6oZTjkCwBCghayeif6m/dw1PMq
RI9n2zBtn67vRWjwm0PTwmsDG8Sk+i5xPl5IHb+BQLHWSzRtPEOOaVr/jgyw3XjrR61ynO2VpHgY
iSJdGWB/GtCeHYu3iVIi4HnlOxKDAfUXSb9OgrpaXhLtilwS9jnpI2hj0x115LvD10W/FjeOsm5G
oThA6gYy3J+bb0U6XKSPEcZWVE7KkyeIa/xn/Dncemgq27QxoOQI78JtDS2vBDsZ4wzxbs/jNJRk
HeyzU39n23Ib9onZmgJHrJ2nYyaeh4fwcRf9vbPHCNQo7BBRQMKek1aztHGmC1rJsaSFgOcQ1sh/
4aJGmDx+n5+X4xcpI8hDaiTFLq0mzRI0n5IhFIiQPSkPwDoSiKDr8aOrmlzFFB9LEsoHl2aa++ei
ObQG/H0pJ4FWXYcY2+mhVmm77B65whhYe5JonyFTuW0bWDN6G8Jxfg6vU2c+5QTrQ9KPxktY6jdW
Nia6zH47IljQtuBY1Rb3V+DRvND6DULaZ5XDp2+sRYc1U0FZS3J8uZ4jjdMn1KgCFzKiMIBXRfo1
4/yhQFCnnvdFbirit6JqE//EC1DEZbeijurrKzAHeZV2lmjHxlUKZYp/IxysWvujqgZu2P0vsMBl
VnsTSvlAnATB1R8XXdK+L0UWNzozwJeU12WkEwE8ccOqrwU6lnFfZ/taz7LfNpwC4E7jklXZEQLn
xAq8lCjRpZboQ7X0Q7e31gX6LffHU5NBQwTnglhF/N9tqCchjfIR8Z5vymIOv4WAWBKbPkG9/uzO
Z0IV9iqseRo0EFxjbhKW0M9MF8fDvFW7CPJJMJCpL+Ljis7fmqLqMZUTqFZPdi8FHMcrX1kdWNz/
pv6Jj+lxoWDP+P6dmMOMTnDDqBjPCqYnKh6k6Ni9ARJNNx+7EDNaHbd4So17PM9Df/PlXvOQaw9d
2/zAuoBuGkehuMrb/mOdsmPV1lWrbHiT4TXFKzd1x8Lay5YunQCpUvwHRtHI1wbqwSPoLWBYjbZA
xvV//GxviEBPBndmo3bFx1wQ4IWH66SG0iHrlwZlNqYY1BXjR0CRT7RdseexmGS9eBGG9SLvtFmx
KgAWIh4zKaCxDAFieGQjNcs3X/2BzY2y8mWi39u2znyXb9cBCU1KzFm07rfN6xcr+Jgo23Jv8jPA
LD1NLyuRuC6T8NCUPXr04yrJ7JM0iNoklGa482YIYHnXMPTRLg/GbmGGhh8sNH1jIpzbngzYQFVO
hTORRoPgK6eFAyxCEtwVMt53Q1XVvQK1PaA90p8IOVBlLgbxwgs2czl0GbDX0w+cqR0/h4Exo0at
y87x7l2JFxEgKX751hLVaxcZQ7F5XDpgq11rwn398IaAlrd8158RzA63iMuQDS78ZXmv7SCy/REw
bovEIay+1shnQPd5CVaWPOBtPFRsDgwQ2kZmpll2ftknl+EvY7nLNDUbXEqhlZ1L8LYIHZwp1Ckd
o/JLh81NoO3IDGOzYhrwEoZ6B1tuxg/uTQ2EH5zEtX41jCYC1TlLtjvJ8OVqziZHUu9/ZPwmvec9
qe0q0DHKUoeqtuZlComPRaPpPwASBrquLfvjWlA4BwwOIIAkAK6kjT7cuL22d2gF9TDq7peazhRz
1fAB0zd+iVWV6NVFi1Yov5jMnYLYJnbXdTomIdpAj2qSeLcjpvUTUfK/50oeKob3Tj7TNLDVM6CC
5GCqd2KM2c5rwIeertyWJBeo5K6u/3k5Kbr8xUi8mgvie9KRXl+7Ht121CK9KUlmWmNh1/acn7sa
wpzEbY45xNRj5VolzotPWQg0pMsLGpZKKkR2pZU+4ZpZ1m3UtmVd8yth4byXzjboq10UAE9ASN8x
jNNcdJaIJsh2pJ/ODSSADeH0uyKsuCcUfiS3WV5pvc5vwYFtCUAhXqG7lPia7ynwsZf0Mp15J0aR
ZFUcByuCs7ZsFsm6I2cOJqP4NZ0AYLvSijNvJUI5B2Z6Ib6uViV2EhtVBFArNxIeHbBUCNWS4qp8
CIQjLo4bY1vm3R36XWxELUZIkX6U6P7MJP1rlbEpD8Z2Dy5aKQ2hP0+BZfSOO7WLOeUizc4ieERA
Z7aWlpxh2Yj4qN3zOdB0z7LbxeZ7in30wc9WhJHeWPBGSBU/301RIKVc9ftwXvhHBiBdaBQBDsvr
Qk7O9OJpTd6w8gxWg54+QS61VtUcCmvV0BusRU54WuQUsnYtuhGttvpK+XdINUhs8g1Uz0VE3M7E
B/UvF2HN5n1SY0N+94rkSAKXf8Htr2HbM+BUY/RVcQ7waEghGnP8Pm8ZOQxavocvVKXabbhHShtC
+VSyV74hxtGfiJ48sgdu4T+q12Xy8yAGD/KYL1f3cNfpi6V98KgQColG4eYsgQ9mcL8dOx9E0PFL
6It1jJ/NaRSeyWO8tAX8BgRC2iuB8t54CJjaTNlVJmvPlqvh+A72h1QdYVpHXPzfl9iAG/XTU8Tq
MCuoKrzWCUxO+bOfAZwy3JHhZJkTqmdPyhR7NiN8frEbPi1ucCfSJF65mpFsTq0+3uLU+E2lT4NV
2jssPP19TfZ395oxw0NeJ6iYwFbsUhuQPg7y9W2A1OyrXZYLSzhGMNROFT30iWNPQYhRDhBveY5i
UXwo7VQm1BU72uAkBHReAhTwqEwFyiR4iG2SbKSHtFxdO5u3vU64eC/JT4u9rmz8pOSvzrTBEhP/
Hv1mgdzsTcWgBB185+iMmJyctbiOOdrYsU5C54qX4ssBDAqroEYyCjIE15Rxamexy40frVmMzwj+
0Dyq3CWZ2CE5l1sfEtT8/MGooBEXmwVbJWHKoIETKlQyF8CydMrHRYCQW1f9D/6K/znzAlSioHGo
DPPmOBO9pukvGBXlTqzW7RMIz75IeK2Y0xxeoZ9SSHP3i7V5bI4/o43YSA9nXZeAnSgUNtlAs/Jt
ZSiGk4QwYIhUtKYth73snh6Mqs4/I20XHXL1YOxV1j8ZDVn7jArGOeyKNu7KLWiLFptOK2EFnXKu
yxs84Wo7dGypGS0fXQFQ7I9bmXVNClsRKzDo3gMgRT35ePOi9wCZMyIP5/IFYUHbKBpN/7LPblNX
kLXUObRRNQSqkSFPmqbBYSsRTJfritbsQHrVgBotQbAX0Q/1Jwi7qLwq/ynmewPpzwg9XuhqfQXd
u/NKgdtjLiqMit9wqUzAmOKTCRseoUiEXASlJAOs1SBiRM/eAjgOsMQKmLqI+AixAbmGIDy0qVWd
sx8A5TeFZHp5IFRzAKh7bPiiNj7lWZdbkf3tyID0INJrZiOZQgiG7reKTcuTivBV+SsDUhGVLiCS
79fXzVJm0Du+6r3d4rpi0DONYD0yc0pepYGZYPU51jo4yUt8cQ2JyliL/OQVWYcXP//XktMWscW6
3J6wdc+NLBgiGW4g96GDqqk6+cKS6q7VtR4Gh9HsPQ690KPDnCXuqDKqGrhQHfUYHKeTBJM2MSYY
pS+Ed9fnuXPZejD9CBPA8FAQuiERwZ34GBf5PRzV9ZLGTKQbrqRTnS4vrZzs3jCVLOWRq44CapZ7
Wq/1uSAzY7q0YzuizU8me+nT01tkFn3ZPSrtx6kx7/eYYQM/GSSiltZ44ba7IRp75ZYhuP9g1fUC
juzRiUM5ETb9+ByhPq7PBzk3Dd4fVX5ozfOKqn6ZuOQoJyVIqHH/YUYe4521JD7D6cUbuBvMkSf0
WZ4oDtWKjjl0u9h8MtAtqqvT4sbedUb0PY84pmrluG4koSSloiZrnlm756eP9amyGt1CNQg+6QL4
awjNoyDF0ZwTJcIahcZAqk5gOC4k6x84FDioMMytjZ96Z7mv5RB7XPR08029N8jnSDBLK43IVHli
jj2Og9+20kuU1oEHTO2mMQNiKL1D2ckIlPNPVZw5oD/K05ks7OVpzYIwz5G894z8OAwvfogasxbR
Qm7ALjUeiUunAO4fbw2hfwUgWcHLk/Z8pzqvAkYXzBd8dcIVr5zwOaRB6yFEDjz/4u6M0JXdVRpo
hj2rRPKb3codTBHfn5w29hvJ648BUbsFsgQfyPLZXdBADZmKnCcsDOKbN66LL/IcQl5VYPf/wd+3
r1W8K05HC52ucsI8IbRCPOEVc+FeBV9aVbdKvM+rLbrDvg7+Jt7kGebyGEmSdcwurn6RpSptlzKs
rodu8OFooIguYD57tRqRvIXVb5Xm4lhfNcju3RR7s1N2qFreUGz5AOqB95ukY7oEG//s0iJhdacf
5pQtaW2ZC436z2FSawL8mmqH5Z5DGWOSN9Qr7orHxqmVeWC8XMb6eOoE3gNhk//1thUZlcHx3rdg
NOT7H2/k6T3zy3d/VJrooCCYownnXtrXWQ+3cohYWF0WYIOteN5xIuJyfaDvyk6350rtdq789Dxp
geY+kw8BInY/FZ/nOAxyG4uFuj7qkwfEnwDDPIcsY+Yask0bY/hIQvoSCkHYuhC2AqGg3va4cpiL
4kP2aSkHWsFHVCnyND92EszTObGBJBzneHvdwJIt7ge6l4+DPfcUQ/jYkFubK/42ISJXg6p6Pl8x
WeTWsW5dopJTt8EQ9IGDRTfmShtHZg5kHCpadMOH+lwK0cHEN5+3+5/U6aHjCkbZdrktkKRLt5Lg
mLBCSyjsd3y5BQgXDF4nelywhrkY4EHeJXhSGvXjbGYntn4xR0+opgT7tuk0lCaCreh9T4ei3c4i
PYiA1gXvwuENJLd+txmrl7ZqynEzcdzJO9VLWDg8niaLrZyqmXG1ueiJaGOYv3pUrGoZEDKYO294
UJf6+v6uZhun8Jas420zfouXEqeYW9A65TuqeHV1PIGyDgs7XuB9tcmiU2LFUAViVAvR3W7erqF8
HvLtTrC0zbQUaL8WKedVl7lWCs0AQI7PCNGcampBVZ2D1Eh1uiSJDChMlllB8ESWpiHN87QOzMkD
hDak/sHZLUWodFdIySNQnzQ9u5KdYc6TqYBbt648xev9aJQ4EVrHOU3ZkGE8hIwMgL+8DveaH2ty
kovEQ5xfW6uTcR5AiFyR2bgs+P4qYvtNNdSECMZhZhB9F5ok8AQRSfxpsnYi2KozqDuB6NbuPitD
fnSNTVKZf6haRLYfnUnRXIyuXWex0o9lxhYQ/29x/MOlyga3hQCuBDG1r+HvLAcV9KZGTyhDn55D
5BXeyFUsEl+iYJYCN8wQZohf9roy2ZkiJhG2bZX4hAhHRkLVHDia7+KP2ty5FXj5VIOkmB9XYtFh
oecvNDkrPjA9xi4UOzQESowcnGYlDYz1j+vO5zpnmEhtYA48aD3lVzlMeg+4/PAH4oP9NtMvg0mk
ZfMsrBAQliSWtn4pgv1SgQRr1cQqfrM1L+co0Qr4RsG7W/biD8AvFELMBj0tAVeHfng4Pw2kcnLH
zgiTAFKLc7w8qyE7vwG0OQAb14LeZkAwCktVvIs5hRMVxoJOaZ9IizNrEcCUbRehaN3H5nq3WCck
DObWpimKoIRBUzkMOLupumTbyt/p5UreFWF1rqU2B242rgt1YfKPf1K/T1zLU/aisOtUVE398ssx
kPZazrgLN36ed7ZCch8EoPJUE0fK79q0MPxWpfStF9UAYst6s/BQZF7d6rLFvGv57Kbs6QXUY5yF
Q/vxz7of1KIqG22cXW8NY2WzsPDo8gDHKM/gAKztzeMff7QJi8jPREWDNB9orV9tD/ll/fp8Yq9l
MfmnOGnKqIy0kOYbPKqok+uA1kAf8BlVVZNzbDAdl43OpwICecFEiz5HSqjYSu1zaf5CBmX8v8QH
aWHbme7EdCQyEj0voMEv6Hym0DRXhO2w5PZHkvCaw7xWPwHU8zH77oW58GOD1aOjHsUSL68eOlQ8
oKvgIJtr3TWL0fNg1gyDJnOl4rsXHLfQRWw4TRdyAb84uOzOQeZ1joVLDCVlLuVZZzWb/jFYlqpl
AhKgM0Ix5yvu9Kg+HLR832KYEQbtyZlE7h+j6FDlflLy5l6jJqV6kFP3PY4gesyMYD1+D2hSyzlU
NROZ8jzAwql19JuOUw0ZZ3RgZ/Xvo5FacEVfRFE0PxGbQDCvq9U0+n2DXNSrcD7vJ5ugzsp8hkq4
qW3fNj0G+8BBFIpPxtX9L8rhy0Fkao/DIwWvWX/fSj6FjrdnCcwF5ZI5E7glpy8zIKi2G6NXbTzu
H5vWx1QMXp8U6i5sDQCzVowv2dmrtXwdb/thdbGOWeEjGQkZ5y4Lq0YhCSgeNuSR+4qv2Kq1P/1g
wd6xe9Jo7M/d+MnpnwPyYK+G4X2eMqvKYhzLrXhw2E5NXn1yqyhtGLmWS89uHsT6p7X/JINBadhk
5+zuGGb5IbV/Ej6xeipLndG0iznTnUIXnByG+4h0xzEJlfuLircPpXDB1wOet/AEr9/DTOmE9WFE
Kmj6Kohd07zs/7BodZYQpOaG7o1o+TYgolq5hyxErAoPr9dWKus1uS5/EPfuk3A+yYszn+UVV0mK
jgTk8B/O8Qrm5aGBQR9FR0YZ1iEe6zir5NfFMMGQvQDlqzlnKo+Rc7YQazaNmMGOl2SLSZxljbBE
qJV8MTpDkeXBCtUMQ4EroUACu0hKV7hbCbHCTLxSj3J6npCLCjegsygj9Ru3s1fWrw9tR6UpdzIK
24gJF458AyKvQnYDxLRiqswFkt/Fvun5fQirhD+dg6bbumcv4ZZTG++Meb5dazXRVQzEI8bkMaWG
pGace5/7WuvRmJ4A8ZutyhosYDCmrVVH+QMISKbeQc60XJIyBhDQ7DYrFyLIBcTh80A2aYzmP+xf
8cgzJgZIlv8Lj4QhBYeaNkWOc4aEMwHIk1CaMqBWV8yrsSYEn7LaUjUwE0zpx06yidTC07GivHLp
1Ip+7IKhzjNSO8duVEnMDQc3iP72kG+aEa7BqxZldObLXFPh/RiwyE5lM8fOyZmPNx1NZAqm3bq4
CsaWkvfUyKpMFoU0aJqqiR6W7fkF7XhZcCNOHgG7IcTLiMnl4RFhYaHaRIwfDk/z9EBeoYMVmhUh
VJ16IEqbGdUuefcBhLUvdrSrNJvCWK9P+DIriEzafYYS3DMKhmZmFJ8pmHo8Ixhqh63kgON0qNgA
QAUqWa5k3caGB4VtV/r0GWeaGTybOKIRLl/7ibQV3SZPSbchF23xLqkX4TyG0pF5tsO4yVCRncff
VLMftTwxj41HPGOLYOfV3/kPU1A9kkGPEIFCcwTqI4qhKaWTyHHRB8uZLIDvpE/dkK3atVF2iWvr
8IxuTQIB8QApwDr3vpX2BlPw/rbJGolpGnc7pmSikxK0yVJ5LD+eblqkW4BGLv8lL04Xsv+6CT4W
lyqnKR1qjFhvmBvB6MfU1n3agr6F2R6sKwNdU0F4puU+IYGBVbTE2xI6dx38m8WbudBBngL9FNQp
vgZIe0zaVpkm0y6kzd7h5hIfg9i4S5zKbQhFfkaG/CYGrJxLdEHKtQXpuQHoIkDHx2XxiPhlqclp
w49sALcBXOWI+RQjr79EDOoVe14KeUzv64XYKKr6YTOMN+Af+kNNC2zCHTbwItwbwAds9Iuu8gPa
6t7vBptejykpccdkqXsJHEF415SGh6B5KNkR2L3ggt4gbFTaYPx2sZmj8j41RG2C5bUNjjkNHanY
ciQpcuEJnCFS1ekydKkhgTWm7OoWg2Y8aXbEQx+ADJ3leXVF8QcGg7lOmKvkhuJVo902ewcaSKHy
bX15Y74265/YDzdK1qR+DUlx5Yqm2FU4BgD0RW1xrIQ24puBe8Nfh3CBirM/E+xx5eHmxCdzHjFn
LFmEioM9Jux5Zx/FdXJ1w9m2gh3bjXnoVKlrZQslgJ3IPxFOAQEYvQD8Hv8adwJ9zMB0Sjw07uAC
2E8q9Vku7l/ElyDAOEmPXxEscFI5/e9mGqn7FuhOauY0VgKT6DynpT6X9O1YhWpHy5CAjOprWvIb
xHlzoWHgkbQvoPlgqdx/4OJAQyEmZEKqIUd9hkSXBhU2SX1be586AirGn5O7ix8oam+VcQMgrO8M
lmJl0o6+3xPvkKL7YzjC3DOJgJ1Ckj5Kslob49Zp+CGZGVyKu6urGGjDdaMr6iFS80KDaFpywhwv
Vns97P1SqxlJQ/GwpaNzfvgjivzupV7YXClcRG0QpVvvRybRtSciI1qAmnL8dcQ3BVvNqJ8gxGGE
Ywh92ZjNP1TGfzxL6jyd4NWroebiZBIO+zi2bKJYXqabbcNAkRDqh8wh32n96ntZWLO5gXW2QXQg
+74EVeX+Mg0EfEaji3KN/BmJotjeDx9Y7etyVCBANFitPfW/IRswBwwtPTTPkDfYL3Wuk8nx6agf
8IrS6jkVn3oNyD713s+n3AkUXN5xJZQlBbryRmXlnAk4idOS2wmyvX+jeD34tAFnQ19WMwkKXxV0
DitcNyrATdFRRzy2IiNjkpX5MZJE+Wo9a0Evr+eNZhwUe5AL0H0wUrZq6WPZsrqalnHvAmamIt8V
KUpw5ntHL9MbBX4+LoXH7JZ+C2sd69lqDKm9UKnFyKrhz/8lZ3HvC9eHxMoTPVk5j9qWpEEsdcwJ
6jpPqUuWeMSD5JTuLvvbprvFpqzOnvSvEnb3SpZPO525AqowBDOf0I5/QRIzytjtXK+ABO5K2YZb
dSYd3JSQ5vN+PonQzvTjUNy2tU+HLQ0D3EliJhQHGl7PJ6pUJDZBHDYZ6El+QByA/S3h5QL+Os6S
b0GQCfdd7dHeod5G86LqaTkcJ2NPFLZqL36ZcPZUKHennCY6SbRS1Seh+OtMkJ3KPHv6tDkVGt2U
n/J0FX82UurN8rgh2Cp7nb0ciNfU3B3br0JcJfS9qJmWa3r179642nIA6WiNr228O9TRZMtjcX7K
dkMVV3b5wyjlOSBZ3wRJkhmZow4sPqR2wOHhSCU1BpamdJ4wKhGW4kNbz6HavdZqFms6UMeK5of7
3oZxLPUOOBICYKNMM1mjLJqRuzZNKXVpW2lrAQXSRRY2+HB4MwxOKFQXweJknM3NpGFoPtmt6Egx
KLnJvwxDcmpe6Lzy1N4YCmZtCyEuptbJAXz65xxvxPIVU8I+Qg0b8iNyp04TN0gBfBlOr9fVImlh
uzSPH2DGRgngx1HeyW8j6OX8GRzw0MW2Cx1AIZpRrzyDM88vjgqRilYYDaYkQqnxsdRC8JBjHwH1
yEhw25LkeOoCabeqvjmgLzXpaqV89gbY
`protect end_protected
