`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JL1bgZMx6U/X68gqWYEktEeyyqogxjU6605fDMFU02lleo6HD4lzSSgVu15+6eh9MhyqgldeM/6o
I0kVXr5V5w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hPwPY8s4HGGCASWdsZM1chsYI5faNryrLywhhOe8pKC9hhGq6HG/BWJNQww4SuZk0SOGqxGAMrRJ
4WJSFCIsCENQYFOhjV9ssmXXTr+yHnioFOYehmB7mvwvpnMjDZrZrsb9Ra9R+BR3JdU11UTX96BB
8huBSBhYVB5X+ilDRs0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IeQJymaodDStiUSbw50TxoTGG7Szf6kBlERO2XRm+tNT8NZIVKGso+psxRlFxY7BnFPBkLwVOEG8
NP1lu+LK0PrSJ+O2LqtZfosASdiWrR0xM+VgOtoOeDTDqe5qjtxywkvFWF3s/B0abwmkjIxJ1uaR
Rhe2AKUUPfVjIrIv9zVMzELYW6VyF1faCEy3hcy02aiI3gcpgky7yPi6Xm52tp24Uy3KfxeZVlvM
6zwO/qjskGYC0OaVImySqBoIJxEFK/8XtO4uNH+a+vM2U5Eoq8JFl+lTiyQYBZHXusDG9VobgswG
I0+06i9HGJkbJICwpb/Wr5wBpL6fPACd5f1LJA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RmnphW7rZitNwqH64cDbydqyt7plkfMs1MDGaRvPU/Y4Z3qrtDPaDvfzJbsnhWlgfIA6utCuyP4Z
DgaLWk0YOv2Hh5wu+b+MLLVczoPdISNQsZSvA27K7x94zv/M8rOFSu6UgG8/R15upO2YLPX4C4ba
cDrKAdphUNUqxMFaKE4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sJVNxeMQSQQ0MXFH9J/fkPXfuQ82wYRh8U7a+6i8xLCVQ+CekGgLXVA2Ykjq7RmYLUK8qPkMEIc2
hI9HRK0lEKa3D4cnrfDD99ZH6pks0XxhapcodJ45obqIffPLYIgrmq77exSHojpKCRCs9dZF06FH
TvjF3b4G3ti1ErrEn/j70YF7SAtkLS0DqSIvatTt80TkiqySMZt7xoXPN6Hb0uuZYvxPo6kMH2c0
vUh0Cy3ZadFLcRlisNPU/USRVXcLmRrLnqm6nUsiLlmK/9LkV/cJI0lvVsLqbfkq5YyTSnnsnaSw
OJJt20lmQkBHtWSbP/8+XNGGWKNXZ+j5C73BGg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yb7swZA1gwJDlXI7MnqffXOljdXnAsnDcaXrwWArffm/68KS+fEVfjNImkcLFeOpU4vmql2e44Jr
i67oTImjWAP01mopJLR3BS5q2jb2v7xFc+AqT6a1NT8ZCs8HHxwVA5VnAtBuEn3CIaLggbVDk99v
IBsvfmnntMUf/Rsf5GeQWn8CRkTV0VaMhLS8H9PozJ/C9azQWK8FoFaNW/PtAQipOZMNUxIICWSu
iS4L55ygPvN0GD9+USVPq7Fz6ek/j8Gjz8PCUs3eUIFs8NQwv8PIQkirpjHhaT191ris0VvkNHjA
NJCoKeKbolTG+bVmJsqBLQ+FPiYA4+Ag80oJ4w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103440)
`protect data_block
fXPhWdjnToRtA8E5S0wjVw6Nt8SnoilON9DSA/d8T8889SA2vEI2UvnmkoaS44GRoAl+/2nX4BJq
MEZgg+CFJaWAQ7aWHWn+WNA9YM0dLSn5PpZ7Rsa2BRu2RIpTIHgSIsBMVJTQpwQvobejJ6q7jFl2
wSdJT9orRQUxt6wcPJsG7T349ctYpXxsy5AFBLLNQTQ6sPPwjagPA2HNldHYRLlrF+TVlVu+6fPq
IkLOvhgmx80nZ8nn4k5Nw8hrSOvLwyLqN5PNAYU1ZoOVHeVPicURf/YLWjrSHaCb96bkioTzvs6h
85Cnyujx0mW391LRg3yEwMkU1UhfkIalUvUNYz/grA1rDJG0zZgjIm5biWtmcW2i+2RsCMVQafc3
jz8rwHpMDTu1LKjoDm6Ui/iZMZmx+aZcWvNeZToMUZ99p/p7IPp39ZoxzY/xwtiEgv9zjlly3Q7U
z1LFwXJF9SblI2khM30mnIOTj7T3J7o3PLwWbve2l+Qu6xa904Ld4M5fNp6LZX+YZMwXnDKh5w+z
i8po6t6V3uaBf0nDVjTX7ALYfa3vR0vsn7r5tw+UuQJCikrq+1solVl7z44CDwujJiaYGykHlPUO
NJGlD41+KG4xPHThOmmuVo6cQmaKdo5xuog7CZTuH44dArN4QPq0RjWbc6CcqC1fU8ZC0F3RuRjI
MmhKJl7BpJH9zuBwT6c3LSDS0czYpVy5l41wMsxA30+T+Q0h22je+ED+4czYa7sx8cl4pjfTnyRZ
cdGVUI0V01GSuUcZyoEXJpCuscaAFQx+sh2J8Jz+gznkChUcmyg4u+wro2wzbWfNQpqp+0jCqlE4
2EkJsCNNlKtuR9Laymoxsn8aKAtHuDzSTMkl21HywGGPCfT1FZdOaMgfrBVYwUstuEK91Z8f6XWZ
ZXuNmFgHecD2D0axpUgP74O1yB0NSTBwuu5Pfq2FMMNUV5ftYWQKAhE+zedx6CsOS44/41arErkR
CxRrovU8EDv/jhSE3dfOZH4D1iC0Wn4y3lxKO60rJG9aTfEeSuOp9rE4dY3HRr1Bkgo2PZ8y4jE/
GGp2XN8NME0dT127T89Xy95yi+Ug47PxG4vV81wSMnni4j0XHrF9gKQzvpB+DFEd4lHVUMUyya8e
Hsk6dLNoYGll0zx1wzM/SlUvyxpdQwF84J7qUPl6CbuwH6GKxEbJRHgBLdZoXVsiCcSmIfQrNrjl
BVL4XcU962gELBa1q+s9caLmoHod6clayQY4f4dfT/jJfODkkJxABiBjWs4KA20slGhwlUD2c0zr
EJT2XkZh/+ciEuAGYMPsGO/S0UGzbbYQCmCJzfMlGKth13OvOC/eMEXKtL6jvZiOLomf9TlhR9Uz
jZrREv1NLIyMWkzWFXEp19R0zLvDpO3/clbPu6pJ3412byTVEUjsBPM3mFiTBhucVgDcpPoWn5o+
OV7iA9uxaEXDM4OkVyD+pLC8lE1MCdU84wd0JGY3mPvSvRT9MA98mm+n8046ddkZ4R5iTKiAcwhk
ZyJFj9aiu+TaAVfqNfhYfCZS8qK1HYGoPTyqVm6PpodLsDu3eQnNDCdtqTSpShPbRO3g+/ABGbUI
/ozyzXX3+lGDsqORH5Mw/W/ze4MDfzDPYc+IwWonF3snSOLLH9/I2ehswpWPNrpT7fGOzYcpoyOh
v6rImGiySU/XZGT5BYiy1876OyUU54iYuvpGHW00WdEb8YM8aQr5uReFXAOlsKlsBjJ575R807ik
seHB6PO9SGsLuXLZZdt6BIJYh4vPePUIpgSslSXcHxe7MPbAipr3Nzxqk1e2nsW2kSIWLSlD+jTu
I4cWEbNkfds9k90sXxL2KzxrH0JVkhJ8kguOxf3/dqvYnQ0WeRWLyw3C/k1bm9h2yrFHqa8QiAow
zv9iq4U9zuq6z1pPjOpgT6/m70MYl+0iU5sVaTcJgHlt4or/DVX83kIxxpjW4T8L7xpwOiDXAz9O
HTnEOo806gKPfeNY5EXuDOAtOlM/xPVfW8SjbzoweLejX56OcKuiBndrGhiPsYmaP0aaBfG0vHJe
8YV81vnbqkieRkLw5QEX6GMdtthazszSP2wbli4Ev2Fcs2KWOk/QhJ+GkFSdN1R5Q31aRae1Z33H
R0JidTiVGOGUBIqsWpX9aRPRZlSvmlT4e/O37KLzuTlS0zpgINu7eSOSrL7sW938eslh2lpbxBQd
5zHKG9OSsyAQ/AYmpEystOx2vePGkyVelqQ/fhVWBIVdHcypfZuogQqFk0KuXXTxiZyP4p69wrPk
NdyECmppupNMNJ+VHGRiRjkOUXcZJ2lQ9LIVagOqtaESjwyfXThqHGQJV2r16xmm+XiJcThSb6c5
UdEfhpkWF8snuZWAjSqnYT/cp1VdqbVpZ9O/cHTH5Vjnil5uKAsO6gJABGhlKxvo5KsWLf8FjdXD
nELzgtFe04E1dwjKafMEpehYOj3E4eVOoVn+CmKnu4cjA05aA6ppUvirxEuqLD1pCiqyxUhEqW4I
35RURnihmIoR253Oh9POOfi3ImhoSU98kqukPTzMPl2EHONxji4avSAZpwIgyy0ipMlF49ObG5NC
xdExxXHO95tmEJrn9KYEjyH+9grSkKXRSonQq1F0UUuCUartDGeNzRdXEOJXLYrQoOyS9gTjefFh
ZGAu5GkeQ3GWjsBU3KXY8sOmCP6XoF4Rq8N3TxRaPCG1Dtb9/A4nQ+CzagbXFxdo9v3zgpoWzv1Z
Dqfno2qwG+dd9pwFvO78cTIy8kXXunyKheglZbLxpBgiOmVbUWoAhwwYqLnGxDMB9FZ6m1OkyBbM
iogcX0Cx5spX4jM95ffjyakT3o1PC3eMneYcRZyE7KwwaIdRy6VWfVoPzD11zJpwUKKAzKpJQ9/H
slMSOCiJQHBNOe7ij/14ff9uhLx6/0BUeuINWRUPGrY9fPPUoJF38yIMW9DRguejCRBqBnXfIJb5
BHa++uk5z0d9qLietTI1kOW/QcHDLDUEb7SHTP9O6xrbA8UrrneTmuz+OB/rm8CvDoo0QrLTewZT
ouB9Wz8zw3rcL7WkE8uaP1z2RGSM0HIQnZ8NLuvTfm5//J9d7pUxyP4illA2MYS2ggPqWkNT1a6Z
oYmf0Y7aDD3wjTBorGiFi9usXdCDvlrSWb4HidSBntblYYfIVvkCjuME0IitQnrWAv6NFCZDinJ2
AqcKR+xq+6CLy1alYKCQVjsZxqXMlcmEf0ukMxoMMxFO0v5J4uI7jL+xZCHgDlwK6dBsAh1Hwucv
unZpMtKL+XT+ntsjQNO9uvBG2jIr593ORBI/opOVctFtPQaaaT4sjsTMaXXi2exiVTK2ORJP1iVe
xbDAKJHR02/wq32AYExMLbHScEU0wvuBu716QwSHhu5kXGKiNaJEKlwoDGcs/XPCwlO9exd1Bzxv
7sAmNtjFyfUyfDlUb1MXH57F3lses7nO/8/xnqqtg4xRv1A3YJybLZ9YwICgF9UTW2SKKEFeY6MA
oCju5TsnrfjaefSHf23xKrayboghcLDbn/buYSwHiJeL7xGa23hjK4QkEDL7o4EBcPvB7RjcuHOk
3BwVwT7WoCUSGN59Ooaf1pccNZeRPuaSgABorcN+t6RyqYBrrhxrgAIyV+4vuziUCzmwsliMwCMN
4B3ufZGhryQ5jxZs++m2vprAFS2WlUdwbQR9sNCjuKHGtq+0nbedR5GX8423YzD+HdGezeUFLgHA
ZjlOT5xH6aNx4p9f6BEUqRALkohIVwZCLhgfq5JzW+ReOS3S9th0t1G5HZeGK/yT2xf8OkENVf/q
A/dwZTXLMYqBIaaz0jmOgCYVI2EsfvZIk1ASCwZrj+2gO6nO7P7aDksqkDHGvxJr9/d5xw4+ojwR
ZNXeQOkJlsMkSV5vTHvmzb7EeN9Nd/An6msHlh4qcsQIKQAMhILZSLkq+PlxOjYUehcd6G6ZzztY
jwxM2tYemT+MAl5qpkAzumKSoKJgdL0xuSgYfQ3RFK/7ZqbO7ygv0b1X9AZs3LYRzgqm9mz639hy
04rlxQ8S/oxZOV2reUvSV9svBkUsFR7eLfHCv7YGpl9DVlfZehk37FVdH2BNT5EcVWy6keuQmX1T
XAxPaWWTEi4vNFC4wGS7ogbpBllCaWKX6E7CA7wQ7PEfFzHEGyaANOsc9t6/IY8FQm4cBAdLWc6g
js88wGMVhfyuUvM3Sy9Yj3K7In1kLkYGdxwmnXtwerAIuHcYLjXU/t3fw/BkAEPvPEauu+WMuoLJ
rJQjM72CDtU1cyyzGpn6m9w3AfGl3aD+zzGgjw7o5d5tkz1+PMTJCa3hbCtd/x+rU1CQ1bhSrK97
IF0/CPnlC4sY5M/ngr8oS9CXGyhLIJGH/mZwkhbMXpCuE3DyDEN4vYIQCDj3Ft1e12yg53uxRkTS
UuzT7F5/fIEDtQ8prwm9WNylRcdthq6kfL1CggJT2NXw/krMijYpo64rFtn+N9ZYG5B6p3OC81GJ
yX71+4JaPZ5HJOylbwUCUs3mbVUyzC/DKC4/cswrqJXTIVm4gFbO5NtZsY7Z81WgYNptcd7emmZV
zL39XNKE0AvLKGJr1LqT8JdFZZThcUBwqvSPZVzR6W29NG1TlkGWyMN0NH35ymiSd9pR7OlpvCN0
qL1mwiUHt7zIcqa+wWEkI9MD2BxvCVbvSfZ+AI5LZD2g89VHa8RLywwDS64GoNNbnWNFns6j/qFx
3XMpkZSkDAMoTOXXO7z4aEwdzza+N2VOabqFfnF7LcNG1CiNH+TcHq+19OXTR5oSw1bv4HxWTKXw
3VTtRwqWqmlWCSsU4hBdyGZfqodwlSE7AxpNImEKWUdiEvqdTPs6VYqS0S0w/JEK7DsR+HPPUKjk
QbZ8ApgmsI/V+sh/wE8j8elidLHYlM2HNdkEcFhswB4KLxzR70drF34SinibCtmEUMTsfgEytGwm
bCqh3LWKhYPNEdSDut5nnzA/BVAWEfFU4+Y+OcEupYYtE4jo58tcj5Y2dOjjS/o++UHuDy0CxcS4
/FCpa1cFUMSz1X0ne2q+rEFgcExEYzTn9Jy1F7BnoMDUMw721nj2oTkwQbLqg3VHDLPWerPk8YeF
ByD8ld6cnYCt1a3snXjW8Gvkyb43fvyaAfjlHRolBKwgjS24EEsx/NpvlbKDNTNZm3wx94alnhEM
H2P/UnL5dn5vx74Wy02oO2oIQ3cxieSOMsnTFLZUUrahogSdxgC81qx7nr+knJRMRNCpmy6DKbBq
nKdwxBWCJDEPkALQWSIA+ARdABcehmHlH33ku3EXFIg7g+hv1NSNT9rsdM0B3eowAf2lxcbMaZoE
PBTdcYbUEBHTUfNT3+j0NXXtX+ENWhRIk3rNRyXk/341dKgvPtFIHfbh3POi3l8j539VcmIhAk1+
LPMiZIuSkl/bqQXzMEp2AHI4paDvMP9Yb3QAQinQMOccfBWT3F7oOlmtOMHt3fGKiPU8JuxwXgUZ
A9smELdsz1a88R/3v4Z1XbntFzXuplfut3UoKDgvmfwnmXHqO4UwIWv4s6686p+00saBykCGV0VR
MJjeDwRXzNTn892IkvBJVvpBa21sM4Jj/Z55j6FMU1dlChv54Npw8ieqSW6QLDp9wAdm6UVeL5y9
r/tCxipCfdwiF2KrJKLfH0IpIHxxcs+92dS4v/+ivwA7SLbpkQrI6u8IDHpDKhlL45aYLnoJr0y/
y5AW+DdXx+oTkOmHBJIZrGRegk3XgQOUGNPa6yf1pwpwcHuMroREx+j71NmxwlRBlo4EqfxlHal+
8b6K2e1UpoIs9+79OozRhAkp2hhtyc4A28fA243guwFsaLnUF0R8MkCYVwlVdXttCZZGXpZ9pCmk
dxXvw1NsS//1uMMJ6wptw0vvJdmpi9opuiz5fLP02jcwks2UpXeAjWO/yozKD79gq90vL+ORedU/
PNu+py0qQvW4fNwRc18x//qvx8MhXHEu6xYvTy6+5ksVS6tQI5tr26fxccT8XTeePRR3Oy5AC3Rr
Vkxr7sDYeckYFBSncq7FV554031EqpY83w2O9cwWEA1CvuFV7J2ARgpFUIpO7y3feMD//VvQ4OWC
aOVK0spz0mFISWyNItrlAGbI3Csxf2WPuoSENoGF1dJhtSF4/j3/4p0nBEiwrcYRPqTtIM+U49Z8
LZLu4qf6AA5hTeT1l2CJXx/QykQgNnDqD4BBC+YRLebd2KaP1AkNAq6cWOUqd4l6OTLD54yZbySr
bFRwbG2nNT4MGTlssHnGbZlgTk1IornNE2K9SZIzS3xHI8vJpbxLKmEN8Mrtp2vNedttg6+HzuOp
TPrglnGGO9uz88SFX0B0QJ5+I5yp/Rxf0cuhALuSfBdALtyCifmJVJ6DFAJtwrBIUjTKuqHVMm5P
QFhHCk6v6V8kFycqF1Ag4z+Z0XCk32tFJgqg6GH3dxtZOuZ5GY10eguO1KuGiyxISBEGlZxkF/Ci
RXLyoJTmLntJ45+5zIgon5m0aQdU9P7R71WdQjPj7tpBb3nwXpm3x1gUjRSM57Fywy5X3KdTLBXI
RtaKwgSESFKOUyS7EG/NUyumPaIu/MSdtjgSi8PapZ0N3XgtAVNzDXTCDcDzZLbHNU1J4H6tX1nG
0uqfC4uWYJPIYb//alkPjae4rtZKbP9reqQcRQ1JF502+naCAHZ82cv5ob8mAXEcR1GDfSHYxdWn
l9b9zAEeLhnG7TsMJ9KZWxbPMpQlX8NsccU9WesOmls6IkoE25Y5gXpvMPUlSmBnlYNFVTsuAkOT
MxotP2vHRAHEztjvJYg/TQlTZEOqud5UIBzhmY//lxPzno+zXdOqKVXA1L6JkxAKEej+EXUJKfMx
xm1flFoxTfPrHe8Vpic66Om4zSEv36xRdlqsnO3JdIxqKSDh1CENIyKvNjlE6wrhR7w+UFFglPMw
d8Y9gCd1VoxUYyLUMdQAmFbTpOzwxaYeZnNGOTZRObIhAWfL62O6JzfcODnJUNgOivByjuiOFC+/
XriOK9jQrxB8IlNtEyGboS9O5EIMsSXDviONYc93NK1VFCydBJSwy68tbjWHG6n5BLfoMZ4YVbo/
zToSKvsS+9ulIwmuMWYAtDDfGEPbwaoz0lK52g4THLsnd7BgSXzRnw0v8AT2drZtOyHPvv4TpPGT
jyPf5DP+gYT03fLG8DWuFIt3uK/OJ5K1cLG+BfH8tmMblbWnwXADSuXnUZevYKbP+RPNSuEjhmdA
wL9YNEdSATAiCDczsaPcRthiFcffk366tn80BrMSdlIXTCc7bfhTslPCSYfkOycfeNsD17zXim9N
6LYgDGpB9sQU/xv4sbgMbA2Ir8ypePgsqggKysXx9PgZQl76X7omZs/HwAPy9SHF5liV0z0+YbYg
erIEbuZ8Kpuz3fWBl2JwmNupOehGhZ19TOUTQ5agHMdKL4WtisaT6Oc7Mt2GF0iPCBUOPKHO7pim
csSUbWEh3D2AZV0u3mBHjGhUh/UdoVBdw9gG4wTNAfd21q4TYQ2Cz1X1fmLIDypJ9GCJmkR6NiT1
sHz8gb73p4xtQR6E7lMzRD/+UyBhjKn4ENB9ZaVl8SMmubfVJokRYcpfhZF07VHloJoMTv7VvNcl
USloYpkojAe7IuXcQJDyOtIkQyKwBR848zieeFAGCk3BYoBdo2O5Qpp1vkfRCRES0YUh08GCpMcc
vwTwtRNlb+WpbclzMXSoPwOPu2oSUJgEvC57Avjh6Wz1FM07b2/oCrxCb/HovWnxGpTjhMNG7wOM
ad8xPkRa41h/9zvSzonNMr+1oHl1NHNrh+c7RxA4mGJbvIlcXn1VxXDwXopqmUNwcXP4khanwyRm
a6qOW0FSG1DzNlS0t3kS6f8afXPJs2cmLKPrCrHs2jTVkXFtn1LfFtRZCH8qU7P987/n0t28a7pE
K70YglUQkxyRWcOo5uSyuQncYjuhzvetKd0z47aH43a9Ej0GELmO201a0Y51v7miZD2T6q4rvGva
J7FYMUl0ZUrLCKkpmXhgiTS4ZAoR/xV55X9nwfq9B1OQsyxgGh9nL+kK//iqs0DsgBzuMGuxnmvt
TNKrFJpfJI0IAn4sTlnrS8P64lNQK93jghDiNK8PaAQhJ+AjIa5pLzuTeTfMZxEADh/bSgZKY/V7
yfw1geH4xxGVtjLeI5L6G7TlRmaOhh++7JK73IJ23xwyarLJWV/1rL34q6WaYqi+R/ZY/yQ4S4dk
QSpFMutDZGGyTjLDnWwOmbJsM2ckSUz1CPjlmqxRNi3h3XBd+Frg99IAQKLa3bAMi0F4T0oC+6Wa
HtCDfB+op3ng3BreHcBBbznFR4lq71TVM4uYfQRhhe19LwtCaZmjdTYtfYb5b71o6lS4PM/41XG6
9A75FH7uxZoufw9LSmfd90T5rks9jPTE4feS5aXsjyntFYwycReZcg9fJkhEk1JB2nUGk4KRw1+s
n6FwD1LnNLA9hv3sSF2VWOdgRHZ0SlcTPDkSw3fSNm3IUTG52NNkSRfujpZ32D0UaHqOJGa4Lzwi
aL9V36YVssilDsM2TSuU7GLxV/dGPnNEmxb51/JMiqzVI9BZdVlVsIR5Ikm0h6FF4dl3YXXyELWc
dNPNpnCM7+uY9T8UzdQCwv1CSbZPochljPxu5bQKAhVypZIj5D5BAEhTgSIsvQhq60fSxuuVKwqE
PHWm7wgyU3b+07dLkECIcxEeEyxOr7siWgHrABw5NvNX/ZiW6w6IalaVa1ai7vJUJvk73eTzJWOc
879/FzWe/2+JnC26HFXFDwBtNoFXAenS8VpxDIpIGHEbxf6djEf0XF0poZezyF70upH7fO2PLB9Y
xswB3lQz7F4WtYq/XwRr6at6TBNmYu+q6n4wZqmgJrrYTcB3ivFu/PrF4IGnNRBJ/VIKepTSvUwN
O8VwvUEeKQtf4lV8HH6jl5yNcw1Vc3y23ZYBc76y4TCX0J+WFZZb/r44CaQ3Yc2ciDcMNI/bvYMe
bA9dnlfPZEVF6jFZBO6TZu+iGVbLRUU08dtEPc0+5yqzH7lH4yLBLYgypHWr6iu+61ct7jJJshiT
ONV/5n5S1+v11faNDxG6rIPW4itZLCBdE9nx0viWdMfwY2Fjn9WaJ4UYdxs7yNKx6Tzq0enT9K6q
zN4jniVuY+m9HzIWaO6YeyONbYkko+rOPSV1qGLgIRkzFlcPPUiveHS3wUYHXjbwatcOABXqKcqr
h9K4nL6lbBJpN5dSBmZvWs0mdhP1KUT2Epb6YKyom+Tf6DRaDSGtN+VkAtONMS250/8j+A6jaesv
hduSAU6KKnWgvuFdCVI2YJZr3sm+xyeWW0szv1WNqc7I6JXF2xh0e6u1rSFKjNU5RzFylbCSk7+O
QfhUW5kWGcFjz73xqiibI3PPuKhOo2LmXsM5/pVGxKkgzgrsoq3K6mnqtHhf3YMNV3FqdF8JHiD7
HlzbQ7SIGVVjlY1o11IE9DI0I6KEaU9mQ0sRLFxzkWASzSWNtooA/SIDeS6yHO/dUorQurzAjt7v
7xzTD6LUGSTpvkoMM99SZFWl0VzLubE7TrqU681ivQq9t/VArynngD0ZxxVDATlTVZ0PfpRznzQE
eEKiqgQO5/MT/rbw5tW/1zU+HX7PPy3Z5cjGgj++IJSAFqFMfpmRzlMXNZlT2MFERrWrgO0yFU4h
iGSlaxbNdmShVHe1wjwggWEYWO8EYHmFzHUUI97Gpu8d3yST560TqtGxq+/X0x+0IuElQb8OYUIc
jXIAdaqflqzaCilWeK343Ds9psOKe3sl0QG6Ps+azRE4EAHnd7d/Ym+E1KLjwW2JLjTc4/gJsqwv
lzY5V/wtc3WjOagmoqdcVAgdoLEJ40qXuUVRyEz/8OLM/3GGyQnkSscY2CtrsW6hF4pPmM4msRcm
RX0MAPSCrydOUgvNYpuEk6j0nWAAENx4A8lp2n+0wid6lkRBw2zdoGDCDf0aNDD4+rLD0jU22LhT
w9dP7WV+posb2rQX3BSJ1atkCdTIzARpWavGE95+AyxNHnf8w9ydc4GprqKnz9dXCR6ar7YcvdLn
8LWKd8cyK8J+/EPhkQVmAxAAobpd2iXhkA9RinlXsb1LjbBsi9uI3p2mDyQUcVXSNUdWtZlcoPpE
jw7WSe/P0ZIVxyZkPCpDn083VYmxhszuKo9xggdp5i0J9/dFv8uK5F4vZJ6OynlKeRR4XBBBYy9M
SLJmUuDuJDkh3vhrcDCA9ss/ZnP9dtXdtsJPwOyYhobUVHQNY90uutPsScPIs1Uf/aAc7lQqUTIT
TfM4QMpMkXKSGmMqD28NQN5o/PjVZd+oUjafAMywOOnLR3kdMbqSAgCeQ1DhmdhGEQt788j5fT00
ukgHDuzAnNJshvv1DRu0nFKRsTIQmB0BZQr/yN/3EBodaejNrHZuFpDL+vGA2tFZP8mc/J0mX+C/
3hyFL8A3gwNWHn61lyN5+lDaGQEOL7EReIsABV6X3qYW4Gt7DdcxiYlJSmW+pqT7D3EZjE9lSL/f
E4Eoqvk+wOr64UqKI89kq6rW7BhafX971loNz9/nqSdCBS4U6AgDES7MNYtjBkZF8k0BXJwjmIAo
GJcSH+ep7e3UrxjjzSAlnoFl2HtIbzrUjpaJz0yuRlGkL5ePr0TuwsNtjVnzDXaq1kJRGp+vvN/n
YHIJkq454uw8RSIqneRR1w2N1NbGbEiryuFOTZ7cdKjDAjz0qc4GRcfrTyuuL9Ym4s8GKhmK5xne
pdJTUo9YnPupV7GosJMtfOGqnU95wgODWhi382hjH2Q6EIZrZo4lrKsvAFfVPrERqZcKZ2j3HSlx
oapAc8hc5WUIKmgbobhghxik7KHkCrRS6JhvpBS7OCXlxXSS8N0IXqiJpSEFRWZeraKwjDVg8C2Q
Tl5yJTUzxcng5zmxn/6tZfaxw4YZUvvw+fZS+xnMsh7MNFOM7vMQ8bezuWbK2Rx7DYxFzIFjhADg
O7swSYGximntxlDmR6E/ZwPlbG0nN6kvegmZsrY9LzUgFot5MIf2JEt6+J3NlmSbauVceOB5HUjY
Akw6Aecs7aTsaV+LrvnqKMLBBhHXcMUQ6OrZTBj69N10YWI5smU/1aSaVaLXLyjY2p5cYCSwLPDQ
qfYT170Kp4RxggeZ8Q06Txf0HPeURmncUpqmqhCy5sM/7YvIZ9NI9qpurW5eUuEXVgPAvxkLAw01
VCLJbqUvP1sGAe+GrDEji9n76PoN/KXGfYtrujLjCFP176D/7n4fCQBSqZ3aFHncLZu1e0R+/cqB
YGdgYxzHjqhTvu8Eb6yoOYpAM83cGgPkO7XZBzDdyyPtrjGP2SnH9/zb7VBSMjOdDEymAngc8LYx
25h4RY42oSOddp7vQkrFJzoWqtVoz335v3o599kGz8/8/NqsHEfRPmMcsYLd9Z7X4AoFasMJx7rI
cVD8XR6M0DevkuHPlz6KHbwQkQOpdSbQS0bWuiJctf2o9ih7MQ3ZFWoU18g3dhWt1dsobCxM2KIm
OVG4CsZcPRFR3f1SZo6w/qmIX60vDotRqJcqf4fUW4HxIhT8hjOeCMwuRwdNHmy2Ns/2MjlvIZCb
F6UYOAKXWZ7P1mtMjYlRBsSHEfLHx849h1Ef7Y7RJBoR0KY5taMrO6EGM0b+l5cB3Vx6LSVewY6S
AYKBvyk4MoT8hTl9bsd0EDNq/v02RWvqu0utdf1hs92JhE5F4UJ4ZRZCQpRDJO11EM8UImcXXS7t
7GWY+usD5EzTWfb9XNHLPA8Ca7nkaiNLm8AyPSFMwyRk6S78K9bttAqBiDF25o5wY05Ws594onda
LyfAHhp4jtqTtpei7JGS5NmT9DCO8rMEXVgP3NYUg6Unhhh8UdiT7CJjQTMMcooRL7KqaXBwXVXj
6HSNddbmHN1/xJdjsq+dr/hkEJwkEYVdRPK0eCacvFbjWFJlYEB+YPCLXCEeHQOvQIHeV8cheVpe
gkYo5wZWn9apCVsiox3//ip/3Cy/lQfEnqsG2+dx9A4woXZo1/3QdtlgWZZNMIUo7CDkjlCP+VE3
8XJ1zQoCs91FxRzCscUOO3pIfuL5u4PpDkqIZqjgI9FTILylUURz1QbIxT2dhenszDLj/jLakaFU
gu/yh8GH2csnNiuGjSJGb+poswuJDYuR5UY3VdVet9Xjzb48X2VJ8EgzdlMHoXzQ9IMby/2uQQkd
trCrjT8UeHupJvBwUu3n1dfR4gkSzoXOq1uetUwvElsEEX5/+lMwsgZ41cz8qFSvoBn0wy1nmXR+
evigmh8GVIQj9ucFjlvaOby1Zv/mMnqO1Log1lt/rrmpg1pJD909v6JpdJQ20cu10YjJWS5OSd48
WXJBNGAouW/azIy0GbBhiICOSty70CBPwFfCJtBg8Da66lvVcoXMtRvn7avP0Q5wvF8eKKPLpf35
+6ynSGLeZwVd8d/nzgqeR608gXNYWhtMq+Qb76hCQniLeDj2E2ytYREWLy6M+S0O5FvcWVF0DCGj
y1v3Ynl4h+wvUCQKEx6cOZhJgMvS3Wewl4MMQUU6qoM3b68UyI6hDkMbGwL+Nbm8h2OsSh4pfyoh
HXBy3RTu3lJnChUTqrry69GQU9KPXptZ5e+8dyJmuE89VNdEbGzgC14ri4rtATJMbCFyCP1lMB/V
DlmLcMZ7JrRV/CqrqDqeeqxZ10fqs1VuFFpi+tSSVKOn+Cw+tO50512ZiGZcPaOWhYFWEp3NB0rX
nHGhrmx8w7g1Tul17ZnzbmxEIgsfg5kx2WPpMh1mXS02Ql/zlMYXOarMkfWkJLrvmbhkZpPj1B1u
q7P2CVtrtR/AkNCzzplUOCBUK1YutszjFhL8yCy2fujzcvk+9L0D+9EBZNZL0BSkW/pbwGcVlUBs
gz/R0VybeYDNhpUvmer73V0P8Pad0qvGnJGUrkBc5ba1Z2Pr8vLTvb0kyZob9YBjLLIyIys5lnpb
ANB/dFaEETthQECiVDHL3XWKK+e4l8UPCQ1ftR46vk9x99Xpv4lPwzsXA3APRYTWgS/CMjQCMRTV
+J+i09LnlDMf2FRv3UpbVY7wzC9Ki+JN9gwcfsqUirPVHVE0HRJ7g69haGvowM+XTiF6QYiDfo5o
C/ZEiuwneLRScQDcAmQ93PPzGCjAF8aCQNWHlqrvFuDUH7eJWEAoZRFcemk7knZ2Oes+Gavyitm/
KxWgOCqeVL3q8UQ7dxvx1mKdJFmy5yiBP26en6VbNZM33z6pVFy4urSc7MlFRwE0/yCgsAp1r91+
Rmmh3G5eqMHeoIVZRlWKGxrBSVnlPMLjsL0r+ko2vLorM3Jpu8mJ/vtUXkTVTgklo0SsclEuSuHz
2UMH11t5snCOc4TujWTo5SFYlAEQOwLC4aYRSyldk48zPszkSJrx0un4qXl1PldjiGI2VQrzAnfm
5xcqisrQf1z1EOS/u7sywWC4qgGZVvPYNP91UAa0SvEYkN1k3JD8+nEAZsJRI5PH7bCZgJAwETgM
j+FmxRg7P/67v9p/s7UVl7rGxJeSlZlZVZHcsliLp5o4c5JLhNoeycuwKl3T8igbLz3+UhFOlNxD
Xlt3n2TJhL2knXeX1e2/WTCzt1lInJuABE4SOVdyXk+zpXVJDdX8YztRp/4OIaboNuPsz7eOCebD
0CHztoDDutHgNUWcsJxB3GK+P39/YtcPfgQ7cvHl0Sm0z2xkAhfY28ACqWHgs30h4MKCvabjNfXY
XBqtR08xe/TWnIARU+kPCUdDaH9E2azxZwE7lT3CXPao0b1z9qGvx0ikWzYuPB+/xd8OAbF1nkFh
Ds3hCXm5CGXo/YHfuM6b3IFuQVqbZkVHC9rYFBQeEFpsIAeN9IWIuZLragG5mQDkTb57k4yKv0Wk
n4nZQy1EegfK6+K1UAkN1R08AGsmETADA7G43oj41URZq7vvQzJ04MB8quLX64hmlrk7xxQl1IEf
l1jbqIYCjpKcLXP1VgWr80QO66O49IcMK3SVTE0MuGn/61LJ7Uj4dlQ+gFWt7g4134BFvhoVGVPD
FXxwwVdhMwqp5hMLXdSBobS5TNDMeVUQ/ny/r+It3KOvshS+D5+PfGGn1ACWDjyCK1UBhaMxWTp5
V58HXVskpANYfy/+lDuIrSb9N5JEYxIHjEO43Rz1E6fZwk7gSStV6eTQIJozinC6hG/xp35HlEOv
qucb3FzxH8EiaZEYRom7gUhx7c9KbPYUH65RNiqu+YwR8pJJcOwe370OwQ3FtFi8K+9lnrlaGtov
mo/eXVjA2FhT9N1/UHcrcSDWvHXcJ6s9x/ZPGG1S+tno2YFirMYhInJRZAb32O4cH74PjK39YgYo
ayv8Grx1Km/pHhSjeSCjwSFV5qoRzZpzLZdTA5mtBka63DmOJbnk3Ox8Wlk3/bPb2zgbDcUiWnCl
TU+/VSU2jm8/co1Ysj7d0GrhcDVRou2lIQEJ1AXTawdb0rb2Rtx9IONQ0Y97h0FIOXAAQBHcwF7t
Cb1RyhwG09ObnfJPKKwe2SG+tMF9MYzY3gz0ojNG//WxJUfdINJFRWacSxKTuGmpkGT0JmbjWecv
4PzDwQB7ShoOl0QLfnvV316EvtafBnznev5THJDmzIDiLbHuzvFo8rYtmManlubGtnQv0+xcY6r7
FhXeSPqavrWBl66w2JUkEU2vyQJp9D4+GE0fZvBtjgUHQ6bMcx8zC3kKSCcTlX1Xc5hRGvaNnfjr
wZOvtCzb7nQczCYB7hQz0qdUYj24heheBc2Cevwb+wI3ZIlIXPRMCXsUoPU90i0nhWpgEKKnsfse
75cUQ3LGlthKzJvPSfhudGm5YWbcnSafhusthHYli4/gjrAEb+bBSyxCdi01MemotQvvuvBMcwBP
wCdxo7OJYtMIrTZPCe/wdQfHHJQDs5NQ5adZKYVVCJuLfdUgCNgnRa5Gwin3QsKNfDJBaUW7Zyxo
7amadPKAecJcS2ZRcZZ3saHfKN+cUYCrQ3EylbRqwD/6welCtpvSkWkpGhBW3v7wlLuPLXxSQFzn
M8yUu4ajd4QUDpkgwTCckWqPQ6PBZNteL8CPT9cdQDCptta1VQu4Lzb/rjx6vwQcagvODPk2sZbd
kC1RT4YlscgCxNQKbMuZ1TGHzISVXElt3JBJhOM455Qmg3VB2m7QGB3C7Bocm4jJKyx58LdtsfiO
PzjX1H+R9CplerMCCtCfpWuf4MYgJKKlP+ZiBcL2Du8zxQIkoOiHeUVWim2c4GOxECeB2VtyJdX1
d1/me+XTbt+uHHytAwSF0vK6v12EJbAtBa2bgBJlnuaLRZQAtmCIyNjV9HXWx3x62F10W52MpdVp
tz4638eMyv0b4bNWI+p3ZVVyDW09KJr7kgiFp1UpW5iEBa+W8va7MIJah9iW6QBghLQheOk3Q9KV
0GqN68Y2b3VQR6YjNwrOlrAtw05I5/qA9PzXwLjDAmFujMGyvbzFAgIQCOHSlKo3VbQOQd3DLMpl
kjXzYN2Wkqt3UGeg+q04fgdoY9ZBjMjajfnEE29tXd7f0p4trE09uGLNmTiu7Zap4x4KM87RtG4n
qnpGIpBhE0RAAy09/UNqtbpiVay4KG0i0mhal9cxGeK1fEwPoFbNEriRKWzuvBop8tqR4vh22KXY
Pr1f/kg0vH5L5pb6rhLfGXW2TnsqPfp2hh/UNeptebCctgJSuJX+tKMoSng9i5ok/llqKMBuI4ax
qjOyDRx1ez4nlzkbrifBw4CcC963CYxXhzVyrEJfIDeYrntXQzywV0nFUEqiYZ5MjwV+r2H70uJu
fQFJ/LELNVMOoUJucrm2j2PvvZvvYQrvGgj0ePA9P05LsCgbN35l3PRwPgfbJyY0NZj9V4QpBd71
Ef9aLD7T70Evm9rAVmFNuUCaE4fwN8oMkbf6PlfazAT+6in8XBgsTdUg+XXtBmusVMxJ0wGlHDbV
jyZt4W01nVdBodeJGjrmu29rViXK0QElUq9wlCNWm+b3ufL1y/9dwwwDogNLG+C+op7olTnhGDgb
MI6EEMbjIwxNBvrdD1OvQDamRYfLl12/TY/nYJ6Ba28tzF0e3e5TWr5CzpT0iVj+HsBNdUGh26yw
gF/JwVZHI8Z2lXC8ONGlXQPeFFaJ+6MshFD9IEzooaS9WDvANjUbEcpaonsImm18CgG2ttYvycHd
g1kXfK8zLPfQKWhbNqM4uKOS2t/vxAjiu10C4juG57mPHwmXL1ZV7twPoNLAf1YuuFkibDKpveBW
6XPDxv7y/Y9WFbYX5u5JOCd1696/mhI7637uSO9SAIbh9qE8Dbzv7TssJ3ycroYcwx+D1a8GjSTn
wwUg8l4zbhY5puLYSuyC7GyDu3KLPwxz0MR0PhkhqwfQHFfizHZnDbtSt54ohjr+J5IHjTmgcU8v
y13rDtm+buhKbWpfYbOE8MiRWDRj602Q2pjesDfM0tTWH8jOlucsbPdk+mcapMVgdzsM/Ntt4S+V
6HyCtF0NxIvTsmKF7tjdjLPDdFpI6obTbqPP+WPUgoGVbTAhi7nj5zUSyHMGvZRu0jujz3iRPytD
QydUvzcAR6eBTgrmIA9lLhQzhjOhYda9KdYoB4/oCXoyk2cPLEAJnJA0e97Fr1eDiclbFsr/JPMV
UMH4Dp7VWXPc5KCMSropthrtIbnIkAcG2ZxF6g9uqhoncTDLWQip28MbnYUOEzwhrs2vxWoCqpYF
o8mfH32Kisa8VCunw0782F0OAsVfcKyhKyKn9LBtF8A16eraTKiRMj4Q4UgruOXE6TpXR7tYj6c4
ih8Bgy+U3uWAcFFQdrIaGsN/RqKBAv3P2skgbjGgIqH/cIRrS6pjz+51Qsd28NqM+X7DOiu9X2tw
Sy13KNW7ORq25DaoKMWwZDVcI3pAfP1yViAKDGLmJyABnj65H2ESISPtMf6VLZS9yQKqz/0tC++W
rhHTsYaCFJMLCFYjK7Nm5kOkhA7HRFATLMh6IoZkyRrmYB+ObadZsTWhPkwPpaBD8dLH6NA8vyMa
OaDFwm9v2dNtZUtKk5jDQZftdPM80Zt7mcUhzD91xxVRPhh4H5OV+iyemRrzurElbXJ1Oe6IoCCU
wL2dldlgSS4MJ8WDKM1yeLj4f3ChHifGNSpCYVR6Rb7KeFXPDe6EOfGFDHMuK85UT1E/YL+A1h1J
PvlrGtM8STa2GUvpqRDozJotmckjZ3Ys1SFPxipevE/iq9nFkUym/VpMUsJ36Xw7ts8SYfcIToQU
YnLa7E0uEQdqBgFMb/sXZGvoLWodkyILbPyX1ZUpvLdMNc4L5eVeom3G50C7htxQL++FQSdJY5gl
p5oQg3GCS14iOIgBq8+dM9nNevy38sudzqL+DJennLhk0QOXb77r9HD4oOUwGKBV6Lkqs5o2/OsW
S/gbken2yMHDBjzrjTLmH0URK7XW4CrDy/PnPnwTACRKpdEGHePOiTbSrzXd5Tc0JEQrP8UMA0u1
R4RU49YhwUD1yq6VMNlXtttmwUP/lzUGCjls8M9IAp6tP4UjqpZKZWoGwyLsi9MnPftGXmKCooE2
yJW+qRHQOHkjmt0GLPeSIGn0YmInWXECgcrad/A/8p+wwW7ka5jB+MzMdTo68FPuiqy9W/wyGoB6
uNwIpvBULYdBVuUviGSj4kceWz+vKQ9lP3rCmaieU4WBu48A8WUpO5SAiUAqAudxRNJjVizrx2S4
W/Td2CmCotmye855NQBa/uDZ7vcRlMn1g6STMF8FXtESH1/k1nmhtK9i7P9PDMeX4z0SRD0vepOB
fRj69AGA9kVZ3Ec9znHpLLiD8f0UKNIRIWdkn9V7rOeah5rmKIhRutev4fJRSTMeRBrVSuEt97dZ
QXYcpbzqxM4kjrjn8BKxeaMJ+ImiaWfE1vISRJ1yDT/lbDeCfAaAHYfa1oiyQicChhVbGtqYVN6Z
VX/gETuR0VQI7a9b1iuxXslER3I4POTZz4fz/AKM2BFQOgrCgIy01Yx0BQLJS10plKlzEcwnvgxt
hySceurOqWmHbfIv3hzpPCpPHo2/Z/NVDaWvjSbsOBTIFaqvvIvwhp1R68rsSx9ZBpogh/+hfUxm
6UNhzbzgPIbIBMwryLDRZbSeicLYhaNmU3O20M0mQ6mrZNf624LOJMZ0w0x8gJedfTpVoJ0M06yo
xKHJdgCx9n0Y4r6T/yRvtzNKPr8oPugi14jX8ZObJ6fqU8CxCLh2l643Kiq2LUUf6emoIPXIIvRP
qLSl7RXXUCzcHE6n+2z9NOfBuZh2y8kr3bpDx0Yo9gBgk92X1zVfwMgxi6cJfqYIvEG/U296vPa9
42IDLOttfQ18AvU0GVll0t2b6DoiujcvQmSqUZR3p20EXjZjIGIyM9LUmpLgeJHwwMw5AZ7AF3qx
dqY7KWMm+WQpShfnJKPN9Y1wO4Y9L7ggpRrkTLCJ1BPnfD4ehw3hgKxBN+JpsehAgtVZXx7Fv5p6
NoG0CCSNLnF6cNbCapSydzpVus717Ibh3+GaCCX0m8uGJV1v3ZTlh8MnHpc7/lVD4ZKPnUNNOCjn
xk2/hKSlX2DDAz3j7Pcqj8/p39o8spvi9IS1KebwSJtLWpjaKhSK064c1hnRhtSqs1DuyUe1diaz
quOEDbh0Y6OKV6VbkmPHETOdalE9c2z6X4MBmlqoP/kVKN30VYebzh3e79QE4cenT23hIkALoWnU
ZdOFCvZRtNfVnRBvSq5CvXMGBp81fidbvmp0eeuUvxKGxDVddSNnKXgBZLdjmzvJc+q+IiFNitVE
zKy+sdA+gyQjjtp0wbCQBSwMMSFDyLChKaktpkzuyb4OJBHuBr3RoLcv8HLwvTujw4SOaBIpSVoA
TFEw1fY58K3xav2ygLEXz2+voxrddQWfBUPwgQ24W9MOtcwGH1SKxUPv4v8D8Q1b9bjOyfrWymms
q3u6g3z5gqMBSO0bwbys3yjliHLwBJjlJBtxjrlBpeiuKs/tvdivvEQ6QAxE5iory6Ar3wdsEo0R
zs/IpyFGGkubjqZeIUf2KZpHAcbvyDkk02RH7ayWadshjA6AQnLHbrTsoESEdL1h1Y9Z5mqjtHuF
/w/heDeCqppmDonifKxc7BY/PFlJ2qIpWO+Z3VuBrzP50TYyFfcoIc/ZixhG24TRcvhZl6T2ioMY
uSt4OAbJ3MCM3gXhsV7uSMT00qtFyQiVTbVuiuoK72YAZTMQ4z7UN1XFN/kb6kZVjxrlRcawlwnU
ydH32XamMVPrhj+nhG/KGe+11FsykxcG7AbzeR+YAzj1xo+RbQ4E5ChHUeeqWni/zuFxTaBL23X0
CKhboQjkZhR6R2ZuknDtoRc3vFGgYYRblf3Rf8asfNzzaf0mzWdjZWBLdZkfzl1RV5O1j5xH6yRt
oTrvKCNyimfNxUuYYowcpHrHHyMwOLAN1lFHiBBK9SsV/IqoAQpnF5FPLwrEaG1Cs2diziwiYBWT
dKGI6zHypHIs5GxHDZNk6D89oaFpI+Q5envYwk+66ckR++Ssscwv4YqSOsLgAi548FUAuhRrn1RC
BVDO5XmIk9Y1yYdn0EJ9NikaWJGLUU6Wk1p4kmjlp1C9AUt0oId/N5PPZ8ZT3AzqISyBafVjT/kU
U1qZ4NkarGGEwGanCTjo+P9ki6pzOfRflBP8hpwXhY3HPH460teKNoRgzP5BBJkiiHuPN7mFgOzM
p9YAa7UxYYqzMC+lUxJE69peQR6xgWsMhZ1jBfeeWJk/jEX7GutUyGcDMmz6Z+aVdt9jBjgeaiXB
np3OYER+jFJvO3Exq1ntbUbvQIzzqKLPimukY8UAE16O0Va2wQtUB6tuARGkxHBibyA8CGUix/Za
GZ7rKpISQxJ4beqRhGEiYK9UNa9BuQmlSPPgeMbi7TqcddB0e8SOpqFNe8HDwtgUIZNwsxoffeY/
7y0MKW/o5BaBOIefacNheAPWPXyeMqPpnLrSs8CU+Hq3J0UkUzxQ1otQGCxrgHInuefYuajWx9p4
IgPNirUw3JfM9rkmsv+Etl7aYurNBKUHqXigUVKRvNMv72rpoAqSNjSrG0bpQD/LRbN+bhI+s+/e
W1DYxTesItyvJw3tBsJpsedDFM85ENj0tBEJeLprmz/LgeZSoxyIwob+1I5QvAG21d9ZHsUW50+l
CDsaSwS/DwUUzwKbsI4Pbt4FPFlgBH+fpAqACyVD+nZWdpoInGIV+wokHrWq25c8/eYp3XRGQjTv
c1yX+YYnRr18X073DuZwArYaVOv0kd9zQF7fnQtK/QRbFgd4K728hFpASGR58xUNFNm5Fy7b2fif
rSCqBEurRHcOJluPXwATECV8g2+R84jR6YAHe+CvPLq6qrpvUUrXpnsbkVFc2xy1ThnsomV7a2M/
UmwUrmROVEjGhD22SolUQgihkzXs6BBFQUV5x8njDWljChjqweNnLOIGkypW+4KW/oMy4mVxpvk2
rO4lZGwE6K8V76VH0RqWTE9q2kFdWR/sXHFZyavhmPtmhrPF7kHBw+bUKeVWjbWvlLxGkNUn+V9C
BCviQVdIUyYDTszFd1EajVsTW9b4v6CNSziK0HkKauzf/VtGayCOXXIXhYX5LqjBneV9HLlDWob1
VEqjTtpoaJPv2zuXDqYW77CMWow5HnTLNk1ymyy5r91N7DHxq6uR2ioNgQwPoXZqocye0Is0jx5m
gdwfyCA9vIQlD0JGrm06iz+rAD80dxRJkaUUwlP/nWI3lQZU95Jq5AKVBeoIuuvJ2U+LNabkuoS2
CJIOZ2VXf9Pp/Wfk/x7nk8sDGNYRMiGqXswSfRkU1JjYlc1tzw3u5E1KvZLMZMmcbQWYKMJWivUk
cp0L9RFL+z1hARLfbhX8Bw0KSVqeo0iG+atlpl/zWDIDlMKumMnhae4Wb9xWOFBrZBeCVlYycj0J
baKwnWJyD04QOAT3nQkhdSOoH+MgbeJNk9N1NdKv9K0F/g7qhDalJuDbw5lGWSlnSINK2U0DUIBR
bN2GLR55C2d7A4ACppRolhziJQdcSsuqjali7zpEHjaqyhhY4XxwMyvCsipyXEugJmtgeVi6Ioyy
VimwD9cwPC27q408B5CAxCUlgk0SfOnx2QjDUDmyLWLxSB4YWDC9Iux6r+r+VpoWwI+pbN1DiKB1
7CDFC+r0oSGGIUU7fGmTs+bP+2Hfpnv8xS2K2zLGw9aKMtve5YlsLsvG4Vm7LjroRE9NeJiS5oEQ
fgC0jTmbxQrnOyI8/MGJZ6NDbmC8tCb5oxjj8vTYeZZiUi5XfF32c1yXdLQT8wRoxHVAxzAHKudU
QHRhMDDfLdjmN79rfg3B6jvRwYN5Tnh0kQnxYfEk+A/NDSfCV7RUVfUMWhG/InfeO3nQ5QWnMWyq
8aY12qqNlaOwjren2HlFEF4QnUkLm83TuQN8nCKXNjWr020cuPdrFaDF6vxL2U9l45unHZa4nkXY
R+7+XBP29/Tb+wWQG4WFsjjMpIjCrlQUWHNQLOp4bvazlJQhTZ7iA3KyQV3h+3GcnjJKjjH8Xx7u
hgYcKWWRRS9KXkNmZ5e2f53I7lgMrcaZt4FUOrfZ0ZkQ+VVK5RYRL8Xq2OatfP5/6DFWgxPO+1FF
omHXoiGB3kwo34Xyk36G+KiKeSiCh2kafL0a8CRrzp2WsAKDj2QdTs/XN8QXch99c9UjbJm239hU
LMvYICYjYI6/h8vpV9B/UHpOidZ0ITIY79LcRJvKj9r2grq0rxNYga8f6qavxSe7P0wySjakRxyV
YAazpNAbj0G4zRWCa8xzYvLKurj9UcdQO65JjLATazqfy5eL77/rCQnO2vTyscmPk34Q/HsuVLI3
+nxTjdWT77Hn7NDRkbeIumyiVq/rEuTAqsSBAEI9aqG5yqPf6TvdpPOT3rvi+HjLVqd1CgI1M2AO
9uMxWrY6tgbzAJ9FXc1c1Zbi5mQ7x44cHGC3eJEls+3HofPVIMq1+7wewzBPtkmqxV2yQZaDegl0
Y2vjzwrs6HVVIOt/G55kmNo267TqEGH2MrCPx0LZAQbGuPruq3Yur4COcripccGVJY/lYw9PZEWP
u3LF7xjeYdXLBbt+lQz9MhN30x7Y8scmVqFbjIdUWcH+sPHj1n2c4qVbxhh2E8wD4kmDuwE+toRC
KJTW8t5XZdcvzzTb20QdJmg9y4zp3exrE7sDlp+mlKnJd0ht0nGlQKNT1jV5PZVcJxnWB28jxpJC
aO7pZDSgCrR7VodO/+3ICywD6ZN4rSA4pZ51nNtT2cky9mRd2UTCM3G+gW4UehkA4oVHQ04JSKPp
5OlfG/1ogjcVv0fTIm3vzXxqdrQlYiAcciD6StewFzifGVCAh1UIKesiHgW7xWkyL1PtA4c8P+Bf
nDoq6maE11FTQk8PikDliKPOkgRuRatZDex/4GPMVOAIvvAWlouZPoYeb9yRMDlsA315PJzOszTO
D3KXGuGSod+mDRyEkZkRvBwg5ooboOwG1jvtAW5Jgn/ZVK9d1l+xIxEidZMHX1fNOhwPCHE27upn
cpSfNJfIRm3nzTGWgRUK1WQeiFVF6HhOkMjvIpXktTOtyQ1HBE2Hths/4Suhror0UclG3J/c4XGK
stF2+JBXprwLMUyk5D6ODK4Sgqx3kQk3myu36EzssD2SSrvSwd+nfdDfAY398OO5DB0SxLq8mI2X
C3b5muZkvsK3XrRwW3uHrInQdiGnsvFeFw6YOZ0xbBOjNBFqcpBR3IxrJfidYuX2mjATyqDAwzXv
uboTSKzaP9cGQHR0I76n9Nt7UdHmndRZPa9aXlFlowYGc84Ws/fm9UGUibw6ByqZNKT+yVRgoKnJ
P7zs1Z13q6nzlPdUsb/KVT1AwN4c8wbjS93dkDnBXmQGt51PCRbgGztfNwLuPfIZjIBtdmTkh3Wn
9D6Zs0jmEdMnf5rGyabUQhD8WRXSD9BcewO+cQhCBA0RCOrO7VYwntA6a49nvZfDUxGPqQ22++Nk
cUdBUaUl8aeqEZHtUQNcGQRxtaKR32ZRVLcqNNmaQFwLf/a3X9Y7y5NOuaE6RpxTGxXS5Jzeu0Qz
q075E/Lei4QAHKpJ7/4eJrlC/FwxE5uDNPcNTh0wr50bT9XNuhjvSd+KfRfX9ArRfwPBYIzwmqru
zqgWA7++4OPqy+4Y5YY/0riVQLrc2ro7imHx+6kXSXoIaZl50xqiiMoUSi2NT5jTcJ84O1pEGj8v
ulh4p3Dxk5wz9v2wMmg4feqvHkI+wTkXCGgHbdwhflTvaDouT2bsOUbQvprSpJxoq7FM1wAfKCKU
Ea/u9GI4t8P7dr/9RjhbGOcYbDh04x0isu/+pniLbC0C8ufOouO3HhWTIkEHhItwpOb0YZVR6xrR
AGHV0op2J4+c1Quu9cHUzrj9daOaU/vhFh2XgGdbjaMdFCpZc2yJSWWGZ2MSw9VWi5R8L4NNUDmh
i2Ww6tG08QWoglwRYaDmBg8UllldPYvhBhxU6w10Mw66JmmoTP5nxryfxhYS+g/n5HwaUGiGxxws
TddlQoxWvL7sy4umxf8156vNNzAEpqS+0D4Jk8EtECtfWgefJY1yrIRbrzdJEtvwWwTUGBGKS3Bc
eX+Cq1RVp+7rguiHrcV5+75C5F6C2IKmUr4rgudFNRDZ8tr/xffNw2MUuH7nrgTWERl0KbnNgLWl
J5Y9/BQhA73nvFZTzF7n4/C8OQWhBlQyRnQH95lAwmcu7SEaTbcS3U6RwXmmGlgFRYssH58IU+B5
pj9224JTUE7rM7M4l89aDAWTsdGug5o/fJ9NhIb+2J2oyZKNSiTI24ImPTq5AnVJ51Jv510/U1Ke
7PWs6CJxB/0haRTD4VW9NSWqHTF0KtOMaGiFRnory1Yi3WDyfBcsrIfOoqE3HRX/SHq6mfcNSeXP
wxBXWgZV9UDzYxoNydzNv4nKtjibzsjnKaWrUtKWbWe6KZhgi/aQs5ini87tTFIxSfEYWGqeVVEP
bzxKONaoz22AMosuhnY6uwLKxLtdCtcOII75ZzXXb3nTk4anFcfKTNjbZXxnlJd/JP9DlGl0hBYA
yOh1yvHAKJpv0M9NM8Ll1lok6dtMuPmyyyS09A+qlTxMYJDXq4gDqyw1lPgelYBP8dxHjkWoCfEY
OkhKPetenX5mNFWPG2091K7KopfLWNukFy55P7wVMUrHb0KKcUyl5t6965f7h86PwTaZu7SJDxwI
MHbt0ISC3pCtkYIgzIHWM1iYb9ugcOuk1mNwHM0z9o/AvjB6uaKdZb9Ksk98Fz92NMlVvP4OB0ZI
IzoNS7p7pDyEad49cwoZb8takRrxQ6ZpiNjDeSOp5PpQG9THmcdGI9oHV9p4mjFUCtntnsdC4Xv0
8+PV5Z4CIrJVVUl5/clCJOH47YjyndUl7oqbXrNhOCsRO05/1RID4cKsz29PTCs5IGE58S9XLdZ3
h89UTq9sQd6OPPS614S12oDFflSPd6b3FYeI04glayJCI7psjjfIpJXA7/WOQ2Rxq41/tlOLi9DY
XTk2ZCg8xwrGgyo92dbpoSNRoBcegeKI8ssxaFxnQkzu/5S7k2oCUhpmtXOj13RmFIo/x03Jy7VS
nOxIPM37wvt8EnCqitZCR71DthOwhiIOxAJTR7MVC5xWyZHAAa20lluFtqhuASNoNIwFmQvRjD5V
O61x7gIQdYLTg6Uu7XrqIxT8BaUC0j7WfsxkL3+QP/i6KSWJaDWh7zxqldsL1ke8sLc8OFGrwJvM
c9FsQhBgGzrKyuVinWgej9LyKh5rl8KZKKt3p87qTggif9CYSIeFJ4fzOxd1WbNpqGG5BV0+gLe1
m1EvMJU/gCYAmG8pF1NTy6QNxp5zD1NZBea2ICoLWJuW8VZTG/5W7ePdvND517OZGANpzpC33/Vy
MLEKkOZ/5UJfOjfzrqbTMQ5RQOo9A8Ps9TzRPe8GiDEbCmVV0+k12ciXsxiZPrPu9NM0s0qHTvPg
t6grMVD+P8yQliswzn112YaLqEmdL5SwrC8l7mdFx+WU8N4fQlBjKMZC90XpmfbxCKbaFEXFqI8p
676GtYCEaX5LzajxyUQI3oFY/04kfwRgTM47CMRETnhYI/ZO4sBL4FQV/0qtV2Kn8ZG2cGBPMzT6
2fOqdOzdml7VJno3KmluF2NYmMbByoiv0tOi3ajON/++zoKCDljxo85IZOSlFXlUj3156bkCyORG
H3cYkSL4Hp6MVv/GF8U0bhgCScvoT9i8UTYn05aaVMCTSYGY9gP6f4BudZLhV/pXNMyuqmvru+9i
53PhgJUX1Y8NGD4+i0OvggOb9IR+DmyFSQvmHXgegDKHeIWQakFV4cR9OXgZ8mDJPp0bnAKdjYau
48xTNCR6JYRjCZGwHB3uBqddRKMDMDLS/2DOc70yLn9XxDV4T0lyquJHsBhisN/yReu8qOKvbugV
2/koUG0axxbdDWAX3r/QNAnj8535ffkXLOWXfoMvsvS2m5ahKYeeLqN+d0p+MWFDHUpVVM/Xg3Ns
qAtMwn/l0Y8YmROYxA3Y6nfLrtQQXUtEcHfdfdwfzvGU1u7CBm3c8aIKUfMBa2qA46SBdIreot9O
QWfG5k8wMWy+BoJyzXRJCSLqQgUNV0KcuI5o4giD4oNU2y+y5NV/vpVpXzgRnMd5So+R1mOhNeQv
X3Eb9ACzMfCIUJK1OimzWttruqgXcuav9FdDDoaiksVMKuHT6GDON0OlTfOluRhqRKIVo484fq1B
TNuRQa4SwE56wjuFAGtVN4B2K9vTTjyh344oTLKyXuFOlAv0TiQ+3WpS9V6U8EXXPOZK29q8grdE
C03kJktQqRwiklXgA0TUNhE4gFZ6p1HIauLtT2rsoKV8vuUIoFqaCa5KjgrImNu3qXqFd2AwbyNm
Yr4yd5LAVFcrQdil7juTDWwT4ygPX9c/1vGmbXNgFFKV/kO0XDgU68b7MlwOOrg5iLyK6ceyHb6g
5W9Wz02ZUSyDWK/hV1FI71Wydk/QOkrTeKMnAQdkTT0pStlDX/6ZxMOMGFaDMFIIFG3R62miHnKJ
jyW7EBlJJuiEIXkFcdOn+WiolP2UDHqxhHiU/htVZhPD6GF5PygXKgDZJbbYuLMhomPioRUwezg5
cyMBPda8x5zwz2uD19T3uhOfrJREMI6CorI0fJa+z/2JKFR5B0fQYB2ns1x7tNiWQWBl/Jgey35C
SIK9RVxIZGB4eIeu3xTDWfU6m/RzVwtG078CtAtFdaopLWyww2qT0bY/Y91Jp4TbYRMUMFAsNLfo
xvqSHtDj+1lB15UMVpeLnwLrQf8/DYwUyL4dOv7rvt8whekjFyqDVyq2q/UljYkc5pu0fV+anPdX
2VnvIPs0nI2EsQb5H/qSJM0uW+BTLc07SUGwiJ5bte3DuMGLeigaQGbFbVeo2011hD34nTAQZjH9
L3+FdfCNAMEcFRvcXWlNIp2BBdyLpL9RrdioTDVB6pBJx1qFUFcA4MwYhAHCWyx/SbN22pxIWdS9
7gzo6SGNXVPJ256iF/PD3iMqaUxP7MRdZFiKRV8x+pu30fPH7CGVVTfJDd0Glph/fciITkWxSU4N
1MhtH0DcLSdx3tdCzoYO4mjgCJOzMVVYIsxejdSUzza8DW/RZPmqpunxnc5QJtR6IB3cg0Eaw8hI
rQ/gqVYNH4V5mZN88NTzfGzCdLMs27XH//AMUGJSBAUc1lswFbkJAubPWK94gRoYjF9v2nsm8D36
sikz7KFjFYdz7WPxOWiop3xLKOfnfA9I1LXNoZzObATno9bmvtaSQyn4i9FlkbWdMOlqAQJrEZDT
552/YRHajtycsCcz98vVoiHf43Lvo2GSQcNfHmHgAfyYbPWqroFyN7eZr73nGOe/NjhDC89SKiAG
6zhkukfZRiN3Kk8BgYR/VKo3spyDX/BKsCWeQeWltC3SoLIJ7kC+3z7Pxq5CcZnQ2+sPlLAuyD8l
m/HjRnZdll1Tigv3+PLShyHBOZrPBBEq7HP4jNUVrmxzbXr/Igq8j34EQyL7LGFU6WMsnQf/nQ0b
tcpydgO3hVtqmIh8olOc/HO7TFAcBvrn93NHZJXwT2FYwETKR9XEVs6z9oXZ2upKjoP4WkZuEo2M
4yI7tc7AQOgQEMFuK9bGiegBrdXgO9xXSUzm+8Sg0bTgZCOn6gkp/aUx748tydgkbeiF+CflfcuI
fP9hK+iBARv6lYyUQZd6bLt0wPIn/xY6BW2BrzhC3nuMp2V6qOXEqbIxahjmzS0ZAevJzF0NEeP6
59o/pkYVIJUVgo76Br9TqshgGpttiHTgxmXmAsumlnHUI2j+8Ub+WrDV5P87VZyDB9hVYpm8nfbC
8oXPhcdsCuoVcQYACKqSs113GXPdk6mSnU8DIugAWmaEB8yAAVOq3oeqMqQEel//67I1KWvgYF9B
d+xLMakzlK0ng/a+nX9Hhe754f1uEbpAkwSMPozT5fwTEijIT8JDoa68RkAc12e0TTvy6oge+3ot
HWVam7JIOiOOo9xlR7qtccSBpxfgj7sAbZNdrgCPPpLn7NTTXHxXUqcX9f4Xex0leVaapwl56r6B
YlTo63ngeGSb5xaz9W9GuemriqAYDWM1teRYV0FGKZWQj4dzVowJJ4DphuplQH006lcuDn4MY7Xw
xXa0M60jSLXjG37dq6f3LtJC5Oq5Kf1f/KFpRny8RzdzkdgcG+p8aBBZYA9AU8vYmgw53BqTZK2x
1jDMltGwahP6vr1YapT6QKVF0XgAlCK4b/JV3AFZrOrfpScfshuJBVeD0VtA695GGS79OQk358Wj
Z0zZHJkKihNX3B/9tc5k6YA+7lDfTdxmpT5UxswErs5beDdlgygdKgnAWPopJzKOZx+RHdEuQlup
r0H9DQO86EbetU+5cssZyRv8XZXDBTmhfZQ77gKJbRmCviFtr8dkfKEiQyAJ48POcOrtNHg6/yk/
jvK/tp/hMTa3sJroztpuUo+oSz+9IyHujA6MFIzreJK+LOQpOP3oT21cvYegBGvo3rdeES5IqocB
qR5lU5Z0WyiUe/CPYpVZWrdLpTWhZYCdpvLTK1PfnDVnR8LS36wgv0h8QrUfHOhni8mSS1j7ctcF
mJpjLtBgXfKKF6CjzBVFB9tDg2VZAuDuuz9dE/Iqo85mCDSlAbOHjhV1aapZGL/U5t/taom3WQMl
xVfSbuZ8Lls1HvogTLfj5e/YyrPlHOoGs+CaYDYueLaMMHNbfnr77rHWdGIWQjY2b5/jCdaWW2WR
vKyMHMDD3YKqSsVLY9pqmyxfwLHNasUhnHPVpwUTxcAQ0j+kGdQI4z+Y3UEk/jaYpTjRy8rahQtV
oSa/4XXTTxn4uZ/B1z76DxfxAN82ZhSoN4PMgO27BpIhVWGL51CfOXh5feAiHIeyov7vSlZht4m3
uPPRB2kqMayWX4JiVwdxzfCwOMrIsjpYNsFbsh8E0wsk2f7UD1WA5HBjYlHOFxAYUCSWiAsFCy/j
CNe7QAgKYxUHDTzf5r+LJWV7hcRkZ9b9FOKnxlaWjSiov/CPAb3rJQcVBJrnaAukEHeugelqu7yS
6AlWDZmw+J+sylwbvrPDzOZFF/otpzTHw8ttHhzKIBzMAsp9xjzITq+6aVrS5GAmpwiPPGGt7k6w
sK6B3nUVUZei/VojFnTQCIcmFBgHOl1B27VTJfA4Zkv4iQLwIZG1hOpmZiTszFdDVL0F8QHTBNi8
7DSOX7bgzc0au3d/fTLxUtbVdNfdhG/QFXQQhCXbBNf0/KGKfIRHuu1YvS6wlrxWil+UsfU/vE88
QAl9exvEbv7L1C2M9KD22Aol51Zw0cDt7GadYKn6yKxGpvbu8Ukwkd83nypF3DU3Swr1hLNW7YHK
Dmul0ZEvmK0VyjXbEnL04mEhcX1GCpQHiDhJEuuEZ79xcWOpws3kL2C5zYaQ2Njyg10f13q8nSyE
6G1XrIr8YXWdAhYGvDs6jlm2z3pTe8m6gmJBqKgXShUHDiQOJjRQGgLNzSeh2jV7yJ+FY/bDFuiY
82RU1AL2ARpua54SR1iUK39x9nAae5SCiOD6gY0h/atZZyKgbKzaruJrMDf65WsIO8So4rDpZw+N
6EWOLfIQICzjR6PeVjH3LIVoOoIikxLtY4MrqMvZsAQ4Cv5yyAFsehz/PrZMe3jfG0XGtg5+4cdm
dfvlXxmHD5moMoVvYGnzVFGC3rEarilev4LIU6/qz37aosPcHcIW/1G2Tf3KK+F/c5eO7ChIX//k
HWwnZCHipXW5WhuqTFLg53FEKBdwP+H3VKXydFQ8af38OWDvUgPi01EEwydI+EM+MDPIZSPzZbqS
KhtCbWp/mlCnd6xgTMlbSu9LfpcDoX2bn+20FgJGVh7oyx0ESSWzPoryHesV/G5zroPWXpCUJp7a
G1gLKxg/3xGGOtSK9sp+qItdWpBd9PKAM04OSDW1dBETJkj7hx20L1p1gPgxGsFeJqQX3DMkYfL4
RBvzGCn/pzm58Oj1nQdOVDPtIkFSsrbymXTNMPbOYl9xJHKjNPmgr9bO8oxvr3mvFKhOEVHUTAId
FVSomYh1Tmdj8p+eKXqG1NekRM/LpoOsYw9dUBZHTuveN56Q0kMobYJ/7sVSA2AOTT/lnnCFA1bQ
/XZXDsZ7IEFGqFjSij1/lLhK4cjaRBkjMTOm8JLB0f+LMWeTxqeIfzkGumVTy0CjAaPkKKyZGcj9
BPaMNz6a16oDjdAqCEtLkyU4aFz5NyEOFH3CQH6ZDaL+XJfZ1eHM0wTSOH/yTVSPYeCXdOUrKv6+
dD/n5tja9Hy8iANCylQqj7386SL9s7p+1ONr21GbGK9h+D6MDy+U1A5Z711a3yJ5Sgqx1euRCFIm
ZyHjqEXyBIglbMOylVUiK+pu0T2LRmK7nAPrI0nPZgqquGMmYK/fKPXkVTetklMQNQwTMLvQmEQz
E78QAPtLZv6ZxDUAmLlpnkw53t6clSBN5eV3qOSvBH5d6bhSTk+/OF4SirvMEp4nkOU0/llxdXYd
IAFlXVcThYXr5yniqFQj9WUhxQkXmHSCiYSAlc/v/lFNwp1ALfjNEJ1QdUtogEsavOTz3npRbsqA
Kc/lxEquc7fiO0gpBNAdTn6VGTkFrXLBFpfmoVMTwmmFE+ou4KBJoN4WPn4otiLshsLisQ7dsbxK
Vttztlh7rN4gZWezhh9t19Ijv/lMMbMuY6JpBVXNvuM4kjcGrQnKhGeu+R86Gj0gZFg0hx+kFohM
fSwbOhCrMFMQkW3FB8g9SIJpcsJIA03DjR3g4zRm32y7XF4GkJhNQg4xxJOhJkDunbt8pU+zSvbA
J8o599QWA+PdI/34MNRO8WZc8xp0gF6iz0v47iiSzO1eWB13bt55bfbSUH8r7UKEVyZK6PNonstb
kl90szIHyaen3UZG/rU7qVJRCxT9TInmarwdjDJeF8AE0VuZ6l7+UGqIO+pWGpSVhgsFdjbSTdQZ
awoPw9LzdsE5JmiZc+Lw+5G4Ifkqp9c9pbvXI6t9HmTYqyuIRjB+6+c4nRjo6jlRPhT4B6XxnnTj
HDbvnESuH1qlrrpi5cgfnhxSyTG7+CXLBI3HT1uMHvRGzwSXhTyq9LKT1iaPcoMYInQ4ubJE1YAY
jjTJpZntyaBxT4KMPjSblHsxJmGE2H/7bIVmPd0LPDron6XzkjCHNFEogy+LUBaJaYHVIbwJ9Lx1
zkyRHQAsshOdqSQboe/TI0bUA4Pj1OFMCPwOZUSk/IiHbLm8OBpDxVOukKwBuQ1+yxrb/pG5n6Ru
bneJY1VzPWqPWiWtBbgqsU7sux39l2AF/b2edsPVSYT2+Q7G6oXHaJIotONha87RQyskIqpLMcph
KaBZlpfwwUuqF2ExHI1pWLJGmwD077dVxc90uJveI+ym5VSpeKRWN/6C1ucRo2ZkC9LnrsKm8UAI
RY1c9D46R91Z1M+TApHEr+pVLbIGW2kOTEhJlqJgCe0RmCBfeGWvb4pTxxTpP2cS8GUXkeuu8rGV
GkyIEah+8j0sjEQIzTK0ICY7ppi8SuEGKoj/ABtKA+Z1hMeUXO4YJ0q7sQ4dMnNLY405uNdDZJmd
KZDaFdU8bkDeBBUKwjNUiWQkRiO3h/ulfLx6zdXlq15IHIwaHYJAQIkAQMKQGHWA/lJcHjKAfa3T
hQjUuW5KUC887l0lU+sen600Jv8jTp4ZfBTeCeVI/OGaz+ac5qMkvssNT66Q4J9Z2QmF6EFtXbA9
agGfD8wmip4RyCmxcTmjb7iY5cGIcM3BuuHjyaBVpjVFqf6rskzmGPM6xONCznmzOrVlZ+I+fldr
40uioubr06gGUg55r9SPrzKbeC6MAdziC5naBu8N9zPF1LObXrXQJXodHQVhy9YCjj9H92lzfjBc
zV8/bsjz/8JjPh35bp70V3K4OPO2rAoSzD5xr7yxHFQGiVsVb+c1nSEefBI0hO6ygbB//avKyu73
9GSq6rsVNXZAaCgk5s7lFbEs2/JC+Sfy9KHby/vJMV51UINopw9/p83u1MoM6BDehP3NRTpY71f0
r4qg+OZhsXhBivcCg4uOmMyofwUSCuv8/35Q47FTYauo08T3nDf54Wj/5jarcmQrheKHrYPNk891
/K0isrpqthJ3XIZmnovM2ya91T1exU/ZwTyxJax8uInn6frn5o/ILtNfr0LRXgYHnAMvaeJ1OBW6
jLXOZCG9ZlOHv0p+b30o3ymOsMgf1b3yu7G9H3VqUGC+AZ5uzbaPrZmq4xwuPFdtqPmUqTqMtxxO
SaNARpABbtX0v1qXtDccI2ATQqb9YF/RUgmyNvSWA+tdrdy9v4/bnCJN9/P881NjaLRTkc8zmFHa
QIiy/WKnKGaQbVP4NLlGUvyXTrLImDYOhbqKfHXlQu4cacNSd4yErhbYoyKwOG6wKxKJ/2mQdO2b
Kj0QjOExlDulHeGJiSg8JsHOjrHqi9CaPEqNcNfavTlEaLCYqMArNVlCPWpT1vJOkKJ4W1v66OJ+
uSNGtHEO06x0wcaXm/pPYmem8Ua9kdrKDolzEkBwkeo7+buHVVUFzfOA1UbUoeqGfa+kyEbw2IAr
5P1djmUo9xmxc5imjaOd6hEUMws95vsbf+8w/OuPSPqj4g5iL8zD/013nEbTBTqyBM81NolTDtY2
65ze9qa2ptb7Ee8DHBa/Oh0c7rhMBDaWeYNYRhAcCsGVBCtikJYPCGNjnQ1Qc+1kivsc813NUU+/
WJXzlBfM85yr7HbVnx1qk+/O60KdFX3jOp7uPN7mrNy53R2Ra6yNsCwZPm2R9/MVTiEt5JGH4cxD
bity2oAP98jZvZFiQBYuWPl1AOhzzc1qg14gULCR8MpuAa7LsqOkwOG5OdJ/pPSsajJ9Y3Fo2q/z
nXc5DO3d9jVM0bQhM6GFE0mhxnKCVSzuGesmyLo5R9t7/p1K30JCjHUB9nriwlStM1Z7G2EXKWCo
dqY/KFCP2VsiGE/DA7PL1pxhwMfCfqytHCfnSmFzR7PYgcyX77GhuAa5x+s56gj1XLFzmdj51k48
8EP470+moCph6NRPpDfJlKKwXCFre5+xTt272xf7coZyBlUH3kg40IbSGpDzniNU4TsiJmqPc/6o
1Un8rfsDryowKNakjA62AYA6CZqqREvE8xa5LqmXr405GI/Bw2eL5RDq1SV8B9cx7/C9DbzzCOb1
zPd7Z74F1S+xa65byI7Jk8/asILR1f2QDuNwDP8+HanHMvvr/dYbvOKwBesbXsA8DIHn7cxqT4ND
ZgsHLxu+QeQFJrKy/c2FHh8ixHauqZyjwyHD7O0sJQhhNfRXmvcGyyW4oMU24O+kHcgmd3hCdsf+
Zc8QRLGrdutwOZUOMdRwVNPA5K1YdbC31HV/ekkYIKSbirFk/Y2b/XYpevcyuhxk2jNG+o91cX6A
AlWza23arDQYlAb/EjkJrxxBgV9PvPijfpgrX54kLY1wPdzcUClJ4aWa/Q0DReseI2jqsYPgh+xb
GFc3fOAGvR993I59RsLJKfYYe5dUV+0B9BQXU1SIt9eNCHvZBwGAYEg28a9GAecL4nyBpTU7ZmgN
fxE1MNOCdON9kq7UufV1oVQZPuLEKuJKm90QjN2kJ4B/FvQ2OVpEg3GEWBEuXPBNT+1hxiFA/pXT
u1o3lBx/z5IkBUaLzI7MDJ1Fcb1GeOJDz+3KFlugpPZG973GULZ5cpSd4Ql/YUmQoMimkoVO/TUk
ckCU4SquH/126EuglCOk+ooq4Lzo2xfmeA0s4MEK3efymyNgeBS8gkwakRxpXvIY5OuahIfzA5Em
9QiLxrg1Gk8qvYnixYJSed5WStb5XQTs5Ys4SJMhf9jGKE+/y4XpMdjHHhbK0KcYlgwAsWelemMh
Hw72qLgKmDD4oLIoFXIjxo1YTxEadJbmKECUH4N1xjP+UvMX0ySdLlGwDy1q9A/feDD2/ikBmcIM
BAbUm4Ga+9fGFq+m+h3ALosdnmsSpiZ0x375+pmuXiT7bFXVKpu5wFj+xXzdw1LGiIhC5t0kAa5M
nP8ji3RYLw45IyFSST1CwlWOw7PzZpW+TxFiw8IyLgb2kC/AQ8P+1F/pZ0gsz4R8k4bw/hG5aAT7
kjAlx0EFum+FOe1QO5gkdjCj+s/apyR/TIP5F6KN1vi/8qDDHVb/b4jEia4w01UwhdGMCAVs5JMQ
XCEfC6e8PDlsPIFGYPkga1bp3cre5GXZrlazZzx39GfHkCDD41Uq/nRU2qcbD4xEmFXp+b7sqkF6
ReDuZkNVa9m0bd/Xmg2oI2pu8Nedc2ByWmPl2LG1TnFgkF7tBBruVeU4xr/y0ZeQ/gjyf3KZKS6X
j6uVInOV6qeAfLO68W+9m35+adj9lvDhMX33PAGTcH6w8Cr6n+Xdm4AuIeNN3MmGewApXYJY342G
1QnoYeXcKGqlsD6eRYPu/FooK4yMY1TWHz0W5UlbyxYbUojZ2QGd9KA1H/ntnE7KwfRFNShZKf6c
JiNixxQyMohNBhvs1A7DymPOT1fhjsvE1xyJwTs+F3iOV2B6aVgNZ85WCDz8V9qXoCCdZBRKb8gn
1skOp5tF3UzbShXjzVWVTzaFl976VTNRLvOp8WfRoM/XeYTYtAgcrQ2/LckGCIqKinD5975QHiIL
xubV0cWFTsmY+pS5Dtysgr17wEg3Qc0guQFLhj79vEK2kOE9viD3M+t5xe7P+DBnhxFh2qan+FjV
KfEMfMjiwTfYA6T+qxQJIhmjRrWGDssy1IFSiRWYn+K0orfzVSyW1EiLCx1gBzuzCcGGCsRMH4KE
4+ZrEDpVliu2ihP0Sc6157qKqyt9wpsK8YnZWD2AjtTt0R9t3EE/bUp1mToA3nyEYJ1vXyTrNu5D
oSaKqZYW3ygHw6CpIVdemD9VGqTe5C73uA+kBaWB1fP+/k74kGZpzxNUOZydQ12TzT/xHv7LM1o+
d080OO+IPfF8AUVyer0DYvJesoYU8VanLCo8uUcUboJS7cKxwpFRENsF6iPQDsl02D2Q8Od673b0
NVmq/33usBV1g2O4tcMDScmwV8TrBHLw67QgMWa6/IHn83f/ix29oFsznP3FCe/JRYo/Fc4sMgGm
mTQLb3mh/zN+4Jn+83iecjWmFNfUCAMQP8jfF1Ck++/NJyXHqIX7BX7jJmoxtMo3LgodKKzxu/wq
AF+XxvURAFH50/L9Fg8cg03pPxyS1CmDPTLDDO8bXqdW7AtmSZE4m38D8bNzM52UvVQS3VMwr43l
ef+Kmbsq5cx50XbyeyxbuLzXJnYWvBznEGOT+8nYRn7GWibGApyRsqJgdJL0CPt7YJiSCNjd4TCM
bUs0tn1DQxqTcKW2tIy0TbaKmmN7TalpyxupVkqWBcyrDueBn+Gw3M1JBKEZ2LAHxu6Cqy8KOHa2
nEbPaslM9urAHiAKcykQHCgiMV3KYjoHPr9PhdUbBBDltW489CC8BNalVZTI6h8nmlstuy3iiglB
vfid6VJ0b5pv5PR/svYOHEYXw6Kkax+lTGVdZ6tf29TOeF8WB8XYfXCIxXUdZBzvNfMAX86hU1bN
VETQPvrdDFlapIc/1tGxnJHRfdrAmf3kNIu7A9vETjjpxV6l4QC3xXqevXq6bfLhZ12kW11gYtxp
GgsnxXohwU9n/tncoC2/sXIfK9VGrlnFvciZrGNdPsyJ70xrZ+iPN4TmDpfLSbETDiz0gn8QVse9
ecuk9RtPuZFqEd4mk283RKzRzA82ERTOillirb4hP4rhXYRP69w8/hw4kZNqN+rlkU3zB+qGkA2D
WpDH7RWkCd4uSMK3VfniHrVlCAypsP70TvlfKhk2rTTUEAHmQBPubdqTGBm/7mm2mN9Pw+lIzRrd
C83dX1uKDV0K2uW3AX/Km2lp9MCItjjZABlvrHMR/kZetga4Y69yl4KGEGyh3Qaw0axJWR5rApJM
0fXkgKoWT27Od5Lw4LcAoGFvOVjfjwF2i+o+LEhNtCrKbeqxrnt1dWctvYqJI4GpKYDcUnBUmRR8
7HIE73KulTVAHlC9UlyY07wq72bMF70X6YEx31XwOUGLEemSwA3bFaSm4HhkHMzVai8TiqEudUk7
aA0PUeugPrTw2KbWkI/DvhQylim3wLprC/RNFixYl2RxUXaP1895GBdyeUSo2zyCEmJeNhvPJ5DN
/AP8d/HIBXRiBZsvbGuRXWF32ORAOAIr27+lBOq0ROTfCAG+fIsu0A1tq/O0iioE2zbmYLgpnpkd
fHph+b6HHnBWlRfOFNxcSCniGGe1gwfo3dhKiNcsi1SCXs2kADnfyXOglgQSsoCRZrrXRe7XtGv1
3XKuqmS6NWq1iaKOU9E3VFf5MXySC+aPbE1733V30cIOO/6RYGpuWw4PQtTsCXMI/JGuQQcAx0Vb
u8C9dxsgwCa1RfEVZx4czKN1fJVR4nenqItqmZiht2EWrFz1cly+PFxven8H3tYP7IWbN5sDtFwL
2Sq9FD0wxdvzue/IIKzYpuepUQDBJMPbOJKhrKZSE/FUvBigZ7+xQGxWOlMMMVv2o049CjR9vq8M
hlMLB/BTyrwUpOLV/KCQKe2MnFIEq21V10hMacUgL7ieTdwco8pzb5F0ZcIFJazp1oUCBMD/2Qlu
lGx/QCrKAVTijS2uUnXDkHmnLYDcGUtrpW56MtT7qKtJIjE6+58TaeMChnhvqG5OWJBWkZtyNuQM
DgZqFSaNTlMLZEXKJptoxM36T7nsnth/55s2Qig3fwOr1bLppTGc9sGYKUbCiTYey9iB4Brf2naX
5ckWgFOP1hZH0NGI1qm1K10LJ9j+bWMDOwli/YHaFOMu7C2EU7d5Luq/lkGPf1PXZvXwgmWKF060
ypCxPEcp+atq0VMf6tN7+8dYfJBuEjaIF2DmQGlOu4Wobgwmbw4BI6DymEYClTlhVf6b1G3/63i5
E9fYA8PzofIIogr+1j6HjeMnSRcERY4/C8n/2DLjtGFu9m+tVmh7d4m5AHVsxOLoV6wQpf15wevC
3g12EA7qUoiUSXfi0wiRLo71p26xTSwWxfi/Ov5/zotho4vl561cDoqi6OcVLwk0f5cs7ilcVcL6
Hg+xYxseKRA9n6y0/IHSdCppm1mOQyeX2hVs+cv/DJD2qpFfKDEvU+ted+DDtlYatq/aSrDCKyAZ
rDDNZ3Nh1nyVsDUkmF3WC0mpIhib7PLixqQmU6flVQkAxJS9hgidRy8dL0/aEk57UW67QEvnQykY
UqW7tgnBjgYx/EXVg+BngNIM9vA6dXaStxG1CfPEnyQaIPMfWm1oMAkWsE46NnkuPHrdIg/Q81DA
Rl+5IptMaDoOKppejNvcUTxacnmHekZkFcFPXH95aLmUW99fnOclxR3g8KbY7dUxGvhYYfIvmX/A
ItHPugBxNhIqmRD4c9GwujmS6tLrGjJGkVTwypLPS5eCQ/ZajeBu0Z/XUArHT583O+U6ZzxItKGr
uyQ3IdIhe1J77Aus31Wifjo7nKm+0xPsls7pWHtiDDnz9X/oNaUc1qCBHgp4+GOuyCi92xmuvqps
iBZ/e5a2QQCUvwMzlZ5m1wrWikpTXsXSQgPwP/XnvvTcimJuFjkV5tpGdxGAXk4G7vVAJvvMFLb8
Eq+dIqlohaLgJ2EGE4tKzXYndEIv6LtGHBzw5Be/cRaNsoDWTmeDH+1ctcq/YLXHCB7kahTDXSaI
HBbAXOm7qvp6xKNifwSe/6kbfVSY9pjHVlX/wA3WiGpnI2DF3phHSx4Rn+h975w6gzIL17kJSuRa
xt1b5MOPjddK44JEvzjzSKM4rLNnCV4ago1BBVX0rOeoGId0AKArRvwDLk8tr/7ZARr7XK0WCPIw
zwe+E6k8muUc+ySGa5H/MihP2kyhkSG7fjKxIP+mv6SdZiInXNUjdhbQBlidBVMGG881XZ4+chsm
RzuMAUI2x1CPNXbYfd5HDW25p72cPWctEUjh50YWlOny0xitGZVayUtda0jPhQn3kujCdgl6tqj3
slJgtehjcEJ4T1e55Gc+6B7glcf4+uDFy6cqRXm/v/3IZZVzaUg867hmGHY1oR0JlVJ7ponn0D+a
+ZZIfWtZpzC0XDZeFJ7KypWpMfW1UveNF4uXztvKDRQ5yeLz8qytAbuN/Ischio7Zi5tL+pgzUwH
JUTfBkpIfup2GSTZJYkDTb9uI3zARXeyx81doDA1C1gMn8/RdNF4Jhp0s40XXtArnsb5jRDUgrjM
GsVVS16Tgv+K/6342YmZdOwufQv5NiYnHV1wY8jTP/Oh5LgjZs00BryeZYwudvyySYurftKWlHHD
cKnvp/fzJrz08ac2W5I3SboyO/TwtZ/r60pOad9lVWSsWNJTtiUppP5JyZWXTub027bjOqrEy44g
ZQRirLEO8BTT4nk7NfdsbGetfje/weBAGgRENc/gFJcoQO040VSw84I3pPMaVW10HOPe0/V+BJQJ
gOGCHboxZnvLYK1n/NYChMIaDHk002Vp02LSvbVHpVut7jYGPdhgWSZ7KWDjhebKyJ7acQqYW/PB
6E4F5qvw7xkZ1C+dpGfvZFevHWulB0dv3TfRdrkVcqnHTftsDP3hXWyPbPeF3jPIxoGi0os0YqJF
GyCqyxVc/7Ax37BT+n71VYBL+dNpjGd18rydej9Qy68vNHeXNTs9KsYDM5rS/b7TwPdA+VUslNVm
2sd2Y5mgOIuIomu6wWQvIrgwoXRl/HeHeD6p8oehe9nu3/ho/9M97aIe5BWlqjip70TciOWNjC0P
S6quXzGWPM1uHuPzMWN6oQM5s+sbtPBwiK//Aw7LE/gezV9mffFiz4ZI7Z7YzCLNaMjDZrCxHodY
8gsNrtUkmYD1jwdMqu6pd8WPfGdqlPwEpBzfWbyYiWBEVcHOkn+W1hILUrAgfRKBtyQZNJka19km
jaKDBJ0pmEClwAVC3UPKjASNR9uZ92fYygGnjGRGlvDCPPtAxzbKwipZCgFDHIr5mMML0WshCn+I
p+f/bsUQOEq3571lfI4oUlP95CSDqraxgb0cn+wGuipkDirmiWHhRr+6HrOxBFpYKQkB8FHXaQVo
JAgaFKtIrLPVbg9tIygz9HeFkGprctwAGFGFugFoF6gxyZgweC2hrmZFXOCGULssnXc+edEHG75w
D1iZaQ/lif8fKbKGl/xSM0oK6/d2E6Sk1+kaik25zmCgLageG7zwfJS8erVu6DKWRgxOy0sn5hsq
5Si0qoLez6OnEiNy8ppFazrF5dPEDVLQzEg5KRSxzHPzFGXUrcD4Y+Q/hlip2oSjistMsVYgSydD
7Kwow6upjTzWoUj781CLOfqQIQceADkXvUGJ8erjOn4a4sY4MyaCWER10j/sn+HALeYGHJRRclyD
+BHcN5o5BzXxmA0ou9xcjSmUkwtoGmNrkOkVT0bKA5gJF8lcAyO4Xbap57KQZee73bv3F9a/bRWi
3K+oYbg8ljX/CdiRqgYtx/Qtb8nxESdLPxyvZzLmY17X7aeIZd7A9WwT0T7+KZFh+kWQjAfx/8Yf
u7l84HY6xpqyIKjwAIScRQW0ttDtMUbTzyMg5j8nkuN1n+XPoxoi2lobf6TebnCAdJWvrFzksIpj
nttIjGk6VXnPTxy5WLdmNa2eJQr56gmYUF/SShbmAGMDpT6lgP/AbGC3kIKRb2eZ5iViwDROaKH3
dNyjkcE4PCPOYUbxUravM0iYcM44TaOyogL02SsSXiux0fFfNnA1GbWeH+39aHeDWlJDM1D4hq+X
mOfN3acaZWYAJ44jK9GhvQjBBInfIAHH7gSNP/zg0F7wZPiIyKUju7EXw5gumhU5nbty7kSEOKye
ubd4pvDBnVfbMM4A/fSF2wDt8mINU+drAszYaTZEGjGb14V1UQpcm+ZIySqfEmS033GZ85/gWsH8
ebFHS/LuAQWqwOV0AiFn5o1dvLXIDrEilAuKajjmPCkXEjysieOAqNzZL1UX16rK34S8HFZoyM8a
s/8DDabC8Jvi15GBKE25XI6+5cDVSwt524gPsutcu3oKiVEnIY4FrQpzvCQmhWQci9SyqdXRu57F
yUhYRHY291WmiochkU8ETXn8LxZF5Gp09S31xN/MT5rh4DQuJAUim00DnnXoRIwDMHZXkzcah6VH
HfJbZnrjORzcXLg1psLvDtSxO9Z2wFoAvZG09dZMzV/WRT/2xmLqalHfSTrqsVJ7OV0rUCHvi2iY
Fr608Em4M0gyR98BpQgnALEyrcsK3P2KrjADH7EW/6v3PE1E/A61XddpXn3TwTwZWbxLzzV0wGdh
4RgTsq9do/7aXFpwHwevFp6wItRiJbrZhZMVdCEZXSPuL4KpUmNp/dGdp9Zt0HaA83sGZMH4uC+d
66+ptwGXpLvTUoLBGoj1IuhllaKQeXziXt6P6QP8E6TMioQf+WRuVMCmvY+weAKIXnaZOqXi6cmo
dgsE1oVg2QVEcwNBIZNoibSdPPlstU5tuK3MLmE8P9CKcQkB84ga58Yh1mZHgWppIhc5znxFL+JR
0c9NaMr2/kf1XZAJewUdG673Go/5Z/eqTs/Ovg64VKG4NLaWx7jlBQpvQAx3ZpTnFRp8kVTyBx7A
WPx53sj6znJwypVDOWcTSjNfRQnqeOJbstSEvFTsgFdlpzwODbOaAg1SlMPSTQJxsFjRvE0FvhkJ
Ww1PUszz2WqlORKhXwnZ2oCsGNeQGIIItcr+1uIXK2tjH1F68KD6WjWlmBjTWDBh61C0VAcwu+Zx
l3udiRWcLZMunzDJvy6CrvEOHNx14C9VkIh5n2npiGVqB3/zZ7fcV1bWxI3ASujN7dmONTsz3A1p
ZQKzhhqT9PBOGFWjGw+bHg0pDroC7HEFYzBgnbfqlcVbRoamgH0drwY/LnhDnxQ5lOYRkz+829bY
lL+vIIhjXP1Ib6p1Iv1qWS3sYsVs2x06ffWFmr++H2TcSU48CjG9Q7a554kAlFPo8qe0WazJWQqp
Q2qp7Sv90L6CWgYavfcAAPp2yhwJkC15OlPW973ZwpGjacP9zDrf5fDRSi63cEN/7jdPQVeeDTJZ
qwr18Pr1Ir65GX/kLvao24LsxRlRsXYVIqP9o7HPz9nTEzLy2cuR4GYqIbBH/wjQkK6DmuKuJWTU
/sxCEHRGEhj+AwHnLf6RW39BGbIgAses32gIjIiN/iiyR+AZliT5eNbt8JviaJuu9B9oaCq9uAq7
wEjD8fwSDLuwB6SWIQP3tzxO30nl9aXnuhHyn/FwTgQcWsFOgN/ZA2Z+h1LgYlQmAhpsYx5BJKXa
RS4qGpKqLkiO9F5kITktXyE/YRrPrgZhSSekdv+vjUuzllOpk6ecF6RNBPLCNKexnFKLHLq8ypt7
r+enlkDenCOynE4zAWJj3mv1VUYuElFp9BQM8TiftLOLGuFWrQ/KPdknOaoKn+CWJ41dtyNT6hjP
bdrd6cSwq3zm2Aasu72bYUotal5mQ05v1sU1NswCQkE6icm/N6mNKXjkM/T+4DEvu7c89TKcsdQc
1mwC9dHZDp/QlwNqDKfu3FnbfiDbEL4uJHFbse9nChj+091CBIIMcmzf6DqWUQMM0SvkexxCzk1G
JwG8hSOWIN0fwTNCLYerH+RyZUS24RGwKyYT0P/sLB08h0WIkaHS4fUqgnnL/5v5kOuxPZLUSBOl
j/HrT1nQFrE9WaJ3R0hoIQq7zxkg3LmbA62HGWv32TLjXzuVGbDbNt2HnNBcM1J5PcsBGSfHgqok
lOzeD8nM2E8gEG2MtPieSYNdJ25WjqMZO0f+UZyZGb3SHIw1Mawdh6oLvAPaq54h7MgJ99ozyxjO
LoxNhKdIawEnapbK2RSzDKAoovm7Fur/BahU2lPV/0uRXuAwWJHN6ejbBGmLselTYcHC3eB20hk/
g1W0lMKP5VjYdHqxfjPvk4nBb4pG0PGSjrgVx04/wdzu+K0QcFj4u75ZABZkAeCRK4F8ihC1yWqj
OYCZQUbM2E/h3+CQ0Dsgn0NpkBXOxRvOedxlyzNh43Ud/BorwJZzuXnQNxTo6zHdh3AaZ4z09hPx
ekv70GL7B6iOjYDnnoEHx8eN0nZbxfsBXXCRZP8Gx4VLzgHVhomjj8WF4WfK2h16JyokrVZZfkol
FtWz9BlR+Uzl9KR/iT2Ah86zxff5MPn8GgH8YYwGVhmdyQhzWL2y8KUdKrGNoaSvOQaD1ENhi35q
MlpXtIAfQZH5G+4z4bUsYWQTbpayS8ANMZe/9mhXupq28InHVqpDacKyzhCmfx0ag87xEegTAhU7
BCL+lGL+5mrZj/skNe1iTh4TkDVd6P78jiwLKj+5LafoFuf34UQU1XpcNavIwar0OAWwkOnkVbrk
QUQrXW88nOUb2jXuPvrqa7zTlHqn4bGDP+1yganZZ05LL0UB6aqJ21Y+XOiRwe/RzWic5YBoZHDt
E44OZ8PCK2VNaK0wZwhH0+odRkhlN2pevWzdtyv18NOpM+luDqvcCh81tyF7XNy7Srh1E+/8nPsX
jI8HGyVQLY0JYSOmV5jaaF6UgL+su9izZXQIktcOU0uY3L+KMeJUGAvYGU5KOpqYuHlV2n/dET0+
OpX5FsrjQJ+EGd3d8UqzOzG5z1CaSNYNKcli1l7L+JQGVTil7QW/HcxYBKhTybrdl5vIc9K8cW9i
VLBMXF7L9eYIC8r7kGVHknJlVkfl8TMUc64NMFh3mbyIKntB2q8+JNCQkUnlAEcUZgXefvGMU2Pz
LsuxvuC/CTh7nLskXmEtACDPptStecEd9Xwn44lcbHhwROSAGnpl1UnbKXwBmfvdIigH9ZVp0gRK
FGEMEm96+VgDDkR/h3dVUOdKkeN3w8xWwZKdg9jVgLQl4zSN602MSt4g/gf1cQU+86JHI7lezYQw
t61EvCuvKODlMrdET31DFfYSGumZzwCYH1KjijR/sIVxCeH1rNWISD/LNPW+HzA+7ekGY9xDcbZD
4cHS3TACcB1AZ6ZNplRNULDOkwzgHxQ6/M6EIjDs6hDkFeFE8qpj+cx685DEuLDnQHDBYj9QGWq+
gVdrUdKC6QGX2BNhEIQDMJDRqAGVqFh/bBhpMwgBbcbCIf7hpSA/gT+1cN5bHdWmiKGyaAu7wrPT
L207STIezAepjGEeVnqSeeaD5zExRSu0HXKcN9YuiUXN1iKQ8lwcEg/yMF9SOlTFQp+IT9dJdzhW
bk6jUROZP9yF4o2FbMtN01F436ROHxz62cBsgI1752+qg/DWVi9qvi/SXT/IaeKF4A8Hn79guMcB
83Z5CqEC6o3Pcsy802ZMlWK0HfgFrsKV9iPDeuoQT6owq3ozB+88tLU4kzQtJPpQ1rHZ+DhzOMQf
hgChvrrg3YiU2CkhZ85/q3xFUk4d03Tjv/pIEjso9qNOhY84aaI7HjdOayPLguHfXpxxtHFYPNl3
dB4k1nkzw3LN3t+eA23ASFvMxyiKTGCUhSBlbylEFymd+cKGoB1AuicMxTswchtUeGmh9kO+f/oy
3RcBBkdxlW4l9t9dhNGygYKz1HxG6UewYwZCrWFrqKE6dCOwDKJG4E40nE6OF1/qmcI0FRhNMIQW
GlVnbJu2fzDHv0gEGr8poFKCBLZPLnKHxL4vFjQ/HLmWY5zEYmab7xJROKy0u5e9rkIpqp8yTnp4
uN756MWnp+vYqTOFZKef/3TQuc30ObRKxMOTNNsyXPXfehylmRoWlyRoOAvuzm0Xm3g/zjbyaAF0
bhAE9YpjA446viwEuCMP5F7Yvzd6czbjHM3c1Rgp48bzz43CVKE9Obj+eOJoP6IChnkiYTU+Cl1j
mK5Mj5pO1dX0UXxOEQQkY8I4GF3En4sozZ4oCpi5oFWe1vZ/UgMUDXMdaQpS3OxXyzs8uQjHd/In
A6BQ5b1HAUYbBpkZRt5oi/7WmFFLSARF3x4e69cSMcakC4YIqF67MDBdcIW2hAqK3dTGCxP9I9Nu
bXrpho95FWIAdZwoN7vx+N0/4gWgrkNnrdCShdB7Y1S7rLq75KTzEVXHOLcOXtcNw1/t4ASq+Th/
IZFGpN3QXG3JT3MGzjYaI5KK1KQmk5QZaWa5ZJ4wL9dkvVwvXuxhFbO7LfnbW20hQrt7zpJ345XY
kyEgWsG+dNNUJDWiOVExPrMFaJ1uc6Hurn+kRiolH18igsOrAtAAK95I/tVVWH5qzSYeeVRi3w5w
VODZ8uA/R5xwF4XNZTqJzZnsNVi8rmR5PvOaia4x3F6bsk7k4skCOZl+KhehyRx1MXZM8UnfG1Ws
RUEgsUITKww1cCjvAM+5Wma0L3n5mQGbo9QTSUYTxUEKvkDgwV926Zy72T4UNGYVeuK/AxNmmNg8
dysqCIb8aML7bE7OlfHdmicoC/dlZlavnZeIafDa/2gs0HPMdxZFNOnHRU/LXtqY7mxbn7BY2g/Y
aBgpJfnCsd841fZR0VqkV/2hBCHcFACO0XIG+ykUq9OzwE6NwdsXQMzt+vdSk11kdviY3solCbFR
4yael9BP8/ihz5msymYOCNR/jTmFYjWd4kcEiw7mqvRDldyItrW9wt4eUtRQ67UUky17PIfZeYRy
wt5TgbBBZWEHqvKnjsg5ZYvcCL48e6BvJ8iXKFOYzrq+CdBzkj8K+wNdwK5/SURg3L9hnp5gblY0
Ig0lyZmifNtKPAoUwivmyka1sctopUrFcUCGJFODT0DfnfyF1aYiHj5N+Y7vdyHF5h00w3lLuNJ+
aoM4mTsklXOxoJ1L7YyrBtAqXjfgBOufqJzYEVC4anHywxL7DQSdSJEizpi5dBjDwtAJIQarusFc
kt4KNkFlefnhpg12qrGRhcw1QxmqcYtL0p3iuhC0fO8+EtVpH+IiyD+Fk+AJe+RdBSfTgsAr69Z1
CvsmdsDrr/9Mupwacy/t6ddxHdG5KAg+yr/D5rOPBqIWfMdoj2nSYAuTvW775irfrbARNkwSa4wT
R+VoZYj2gSsK1Ck1nt9SlikuFSRft+xWGAWX7vA6ek9/B4bsKTiBHnv91Kik47t4i1LXQVwJsSNi
6DVt8+2xTGoDE6864eTw/WkCMdBodH8P3KK8pCsxwnRGxNQqEVMWcXNkZRHAOjRD1r+d2kYoK6L9
BGUAHRpI+DHs/6Oq40gCV9azu59OL29WUGd469cacNatg/Uq+vZgk/9XqHYy1q3B7kuLyyckRIeR
BlAAZMo/MuSFA1982EIZuUjsc2WfpiIBLcaKyMqXdWCzoeli+HA+Va+3TnbwoCNVqPvcxEL0CgLZ
cevg+lgLvNTxG3motDK8JWDM8Qt5zu4cTDgBJJvJB51FU2Klr5c/ieIbRkqlHqBwjlsnVdDHo84k
8JB5WTjjLccuE8AQCfFTe5YhY49uQuzxuYsvgcOA/0R9LNIMpS7xwWfwWSWt8oLSzJ4Qk+XOg8wM
dfeq/Qe2iqUvBazGVksNs9N4hSPTDAue3yZJp0dS5VV7H1PGOvVtS0NCtwtW5PX7+R608RM9vHdh
PK84fFtbgIvovKLwhQWp0F2IpFAo3rZW2girftgDmXWYZeTYZFPmwIdSrBVw0rrryDGlnqWch2fq
Or5uLnnkR+zqEaQ5fB0Nym1ggeSAhfhntM+ffY8r8/twBiy2Ti5O72hTCyS0Ng9c1orxUBzmyv33
1Se3NS/00nZ2UA5ldPkjtHgmPHOd231csbXlTi+YNBlumkiJzOULO0zpsxdjWBGAr6eWRz4o3f1S
bJp1mMh1TjJlaiHubrMme9VZU8TuXHvggHuTqvW+bFcPIysQ2wv/+wzOyd7LId9HK6+vlLgmNPlx
bkRTmWlm9/WxFx9GY0ynPIwDB6sKnreSeViLqGi+JBX9e4kanfbhO2m8SvJHlAKSsNNCvV/1c9sK
s4Xjt++CMc5hrKDyyiTb6mE76i19pJTXToaetKpD/hLvloL1XRxI7aMqEQ88dhgWMcBtlofrzxz8
Fy+bLDWz+HIHNDHvsjwS8zwP7moBJ0OmQqcmuNpK/5Z90SI9bt13zTxrklfNqkjdB+r/eul4+sCC
hDFLzchaSu6p202DJ6oraxV1bea76L2f00MfpV88fc0HxpNYg54u/pg3p/Woqn5zS9z+ORXLgLNy
L8/jHbYWg/6jqm7yeDp/s3Go884bqoZl2A4Rv5MqHhwlX73gm8uBDseUZ30dyzg3GYO6HhfjpgGL
HtmRd7A8Jh03HFo50YLmPkpI9kQhnL32dGklzMqIPAigpGyPGB+ihCAgyNrYtxGIMRl8iSHw8P/k
inFpTWWmIJasLlBvf6bzSfAzQrQtRAC5W3qrfw+R+zzQxP+7XVClCB/NAGoTcBYUtafIJwsAOKrA
Ob82ycDeR2XOduxyIn3gKoh5JNhmcfXi6JQIoc900lxDg0mxrL5z9uuHKnMxMDWgHTUzvhuTAPv9
URwdxtU8Eb026hkoL6dt+BGAxxEg5KJecYipX85DnFvlVyeiwJpemNNSSklHb91pDNX7E99vCUfX
oWfkxz0sWDOIpq4QZ+P1piwUBnMvD0wLXvN+kzmJl+Gb8PTiVWZgbM1gVzmIq6QY+sNFGfat6wjV
iFNNrEk6EmYMGxtqDJyDSA2p4RqbHvp8gdxiIeWLg+niWmZoj6g6NiMk4OomqKTVeq0w4fS0a9V2
aLMxIMBPN4PIgZ4h04r9kY6PwOHhchOXHj8N+mLRha8wDnlhgJ6t7/nOD8G+NjeJsLdkQga886qo
TQtfXaES/4h1izp6BsZgj2fTfwwxvOC2izOqPq3OvTcYb0SXoOV4LSM4pwHFBuAZJc7CSLhAnxzB
870NB/dgyjgA/Xm0xmGy8bwVncIgoTcqwccBM/gWtpDs6ZraJLK+mxcQR1o78bhM3n0Uf1k/4B2U
izyd2m69ndC8+IXVq2maw2Xe3j7H837/xYgASVHqNpJuGWExBpf/9qSxKe5SADYhw87OXnYfcXSk
ef/lGI2ZhPwjivTzZSaAroGhE4Glm783G7VAzCs6FM2s9WsMkZbFQ1oxSh+RJwpgqubnh2KLYvCM
slb4WoXdD2tq5v8GxsEqIGCijGLDGamCsPBd4yvB0Gz9rTcUK2hjdwJAjyaU9RV7bC/BSjx8CR3u
zOWoFuHYFDVgLxfY0sqZUgPp9x5qrfXyJQ1Sn8iHomQK7AZssyEx+vJsbVQHsVNlk+O/Rxemx9Y1
qDefIFOa35WLHFvaAISlSMyQby7+z/97R6BCN3ArJtd5PHdkoHLLiprRmlsrDkugi2AD+vTjaD/W
StIUggh9noUgmojUYwBx2nGF8Tq+mDgj+KszyB+h0fnuDFI838iJ0PbpQCBaPcSCe7BasSMzi5xc
N8ImI6RJHHXrH0wPB/UHiV0NQzmIGeRmgfqWDKo0Zc5sQcrUTnp92Fkbk2DVQOGd83EG30jj5v0O
Qv0ekqngD8lpks/vfBbwirkZ7a/Z1P3bQHKa4DtqzFAR/UDP8Av0TwZqQdMqTNVNadlqmkIvbnzq
S5oAgdJ7PIiMx0jDv553HuRv6zrHKtHYLubhTPPBkXX4G43iUXrJ9Zn14+sgPPpbDyOinE3J4FBN
hLjJksf1WS2GZ1PCQH+jm+vr4XuBNiBdK0zdSY9YJX2NPG5FCAJ+TtMVils1TDZBldc6j/QsF7Py
cswXoNzWMIWCd9UPl+gtXoKzzLS11m2PSf3IPb66H8JMOL4WtGM+9XGjIWlNTuozzY+do72mNG/Y
x7O/mnIjYfj155V540rvuDYf5204LUPMqzwMZWGx45dGioVFn7YjT0/7Xy7MYRjMJDJYCMeRIdU+
20dmv7dxOUP2KhZ6YF387VCM7LECzDVisTOb2Et3/z3RBOltzsi74C00TQvTimLHrNV+3AOgB7n9
4B6B6JzlGv9TUN4N+FQ+vhYa0KQKT+z7e0phkiY6EKpcenTWngxsxq0AvU2MK049dm3ENLN95skr
NlTOGJxHNxP6xllELm+hyxFHUHHJEDrFFQFgJUR5piOY7G1gW/voqz1dCSDX+H4ROjrVLbftKRFy
5ELP4DsX88zGnw+9pKiA8zbAbJpcb5Pn0XZAlIBQqdq3Srktlfm3JAYwWB26LTNa5pjauTVHIB08
ofEvEdR1K+oEwV5j/DktHli4AHsIzFhtHr+YSmpnN3VDv14vRYet7JnQgZeXgCAtzu9ZXmuuJ3RG
m87hOOZdZRV1lhJ39NllAJ8Q89h+o87gO15sRbQS9Kyl2wI95aSsdqXv3wycHBtP2YFOmnryutV2
D4UlU0GR53Qd5K3WTcJDe+Hzu67Ho2tA3vafKpmnaM0z38rt0oQIqpJleUQ8XN878cuBthrP7PJJ
ksec6wpOwCHm/FzMFhxD1Ggx8deegO9VNcMEXhudgiSLcYfOK0uoRiZJPOki5EZthTkwe+IpFNVm
1NzkGtOzyEmtwnMHaFMsJtIMJdsyhxDEzzsa+COkxV6oXXqxjMb5+Xw3E5o3xd5o/bgPG1gLMaqB
cXwKZfMBDPosaLUJBISWfj+KXVsZIXVVmEr10IrQqQ+lXhWDbTLG7SPGWAyz3IEoON3w5/jw4L73
QqzBrG1zwCLoVsmxU9ifiyV0q6GZbZ8fX2/iE4Ch3msPsM8HtCIMtsgDknTspeAubaZzkd+Hm3nR
uY4YDLVIh8tYwKBQbON/8wn8H1dQvWEmWN9WwhwGH0A89VviUHAS+2gUE37aLIktB/xWT91b61gz
9uQuhLCai4RSTYPu2vvmK599iLBsNrrUedLN/XCjDgC/os2GKBuiOjeuW9IYthJ2fPN5ej3kkUcT
Y9DT1uxl/9vlrWrKP7PkQ52uupJanh3ClS/P/7ukAGKMVcnRAkvWn15QM4mlwFe3rJW5NoMmiCZs
jtw3iJWIwUFpEMcrfSfnJvreMV/djsyOEqzWPVU/K7HmOfcYX+2g6TmmLr8j+p3F9QraSN2N+84g
6IIouIjzNAdrQ0trzXVWVxjGBvZC8qjybkh3/zqCLUlCrLpag6hZDbdJlTRZsd1Qd45hK4MRJ1aV
u+L7LopQpqN64wDPcklXBrb8tUJR+GUN/z1KC9CwXCYHubyM0/cxWD19yoQzXKRF9mvk1thbQ03g
waq/NRH7Q4E5MR6ENdNed5/qP883XisO0pDLatx02+p9wpmML69jlIbe4ladC7LeTmf3UaBjSNuJ
1GqbqmcO/E/th/JJFWDqbUqHcxpWDK06L8kf6PYHmPNiCD9vAvROvNq1Q+fMIU0p7w1KTgVweTNn
L8vcwbllhkYw2dHWGwNRYc2mGz3h103p9efkFrF71eKOpkmgUMpa4g86+cHKHmqb08tpKcVgQq45
m0D0rXWfZAPhUbId2/4P6r0Z5PGITWg6zp+MuoyYe2t8CRy4a9ZP5jcHUn0OipmEW6ECsB97jCFN
86X4xaFwsOYIXta4b9FHQ2H0h4ALsQCBCgVGzgJW3XcLFlNj+AfRh27RK8iWFamjD46dx0iHXpGA
vhYR4LthzpdtzuQDkXnmD5UsPI424M15xugd2xxTvjO7Gv8VJm7ANSNuICf61fhJICUvcJdeXhp5
PLgtIrsT3FsBLYCl879x5Yey9qbkRUKR08+Z4Rzb1g9Q4EnV0svb3R09odpE7Hgf1icAOa5YwlUO
zbMszjVv4hPhccP0XrYE6nYlF0y2c+q6PPVNeuLnX9yG7FI+bEu77hGsbMNZPXYOLj4RrwwuyVkk
Dtadoc7lqa72RKgjuVRIz3+ApfpvHJ/FK9JuHbmiuLdqGY97RMGQWC97v/qd5sUneS5Ek0K0fIhX
276Wiys0/8vxT71lX2dh5ezHWp+alrqgezhoyzq+B3njK3YTQcfcqIH9FDLdUBqsQKA/Z4SewMdl
4pXxK8KSifePW8SFa+UgQZhj2zQU7IzHdOVY+2/aOrHxT7wlispVVKwnb1qFgEOXZ5UFtUe1bcgJ
qdZpQhB6+fptzM+LqbAA1FLZmcrBIZS3xnMA3fMsYh69oD6NdygiolkNKSmaDjQAbe4aO1DMpOx/
UIYolKK7LrsSfy3gQEn1Bmj0v8rIrpKwifnCRPIl95sI2oC4NVdQcF6Hxx6CPnydGEMjR9BuS5ak
49gsfJMUnyNtV6fB0D8cho1LZ6VSt4QxEIdQLaE2pqnjHU0lFvpWHLd5Ms1CILGqA5lkNHg1LBX7
mPdJj4hpKXFLkjLjKnFdUKragky1F5Md1OTMpvKoI9C9jxrGukimpyJ12EHUsWp1kHFo8Ys5CEVo
V8+Hjhx3fPJGPgiT5f6r8D43YNW9gZCqEMxPr9p3LkOMVbmPJCzMXOS28vN/KkMEZHqOKRR9anz+
Bo1NZklrhjpzYEMkXRL2VjavQI85WgW41WMJRuKtnsxVuDqNi4BlVn7xfO/EwpfjbhDNdA/v8MtG
u4smFd6KuXv8+GTl1E66qZhy8Pe+tXcZwfAPfVM6+n0uwMCGPHGqJQcs5fVnNBYtlUyBRd9B2/hg
HH+C3WjZnvfpZDdN0Pni9UW4qXcD/KPlPbHE707O3Wr3EPJebv4fXA2gEA9R1Gj9jWGH/jKmIQfi
mYx9IuNSMUH/vBod+T+gxXOV4H4f+/hxEiPhaNXxRmOvei4OSwDjEMRPkA7qQP/d3/jgDVmzXTjv
GVVgPY/XC4ohMeTmLqC6KJu/LsnsETx3MWqpd41WDlkXQbcmvd7sorIYnWFtW+C7RoqzryZopCzl
pbuDui/CmSN/oH7CPMfitBDS2XdJm6sx8rWiX3f+bbhBifJ3p4bw6XcK2Mkgwt0RM61D9viwJDLu
FOCvqyaQwgKv4nixGxmJJOKoE0I+v8aHn1lrVWifkANHM2iGfuEm7GC5NwXB2fPCc+GBq1WYUSt8
i3oT5v87MlakCA5roz+cN08JQBXsgFoCF3The/C86dT8jNq2DeHuGgIo0/uDVBaoFWJgy1RLBWmG
awo8++bkuTW9YmF5Wvyz8PwQUY7u82yTvubxSm/EaIW5vDrZF79cq1ai6dCygbC3DE9Mp5X/pZMY
7mh5EdIxR77nteGO02yR1Lc21yrRSuDtXLGBWccEdc91QrXMQrwXExoUTQYebCYKo3f3G77aZ9Ft
DdVEbX7mraJN6/IastHjcTD5GNhXY4Q7LqiImB94Qm8dvaERXQ8vtkunPnLHzVLnaFyp3v8qmqjg
FeYNswsBS382Uga7W/qZf9AU7VbEennwTx7GANkULJy2xyQ/8e9etDv8VhRnMlUR/tGHxmvky4L8
q8WF+JdBM5lfPr6UEqUAbQSHo91Fn7Ge4NPb3Xa40pgsiH9RGmKkqYWOo5lSbQoYv2RFKRjJzmIb
/dAEI6d/gVK2PQ3I0bcbRWvfXgReEVRaI1EAVgSp06zK6FIQjMOO2x6fYGYW8ywDszOvKng3JXU4
45WdF8/DSc174RB7ZocQCZTmseY+Z0gFHR0KarKwj2hlkz0NPfjBtu6vuqjOfaBMBKIWpTj60UqB
CEMLWwa/hfd7upho0bEfxr/Rb7Y5FF1djwpHHC/Lk3zIjRFMF/F+26i7A9dlWMn4mTDUHMJwLo3r
jowWWV9ZjsoHgc/hUVKQehY5Vo4/iv1DQDtPUfHkPe10EqV/rpiShyj0We8FWdJkMkpmijRkGhcR
J14Ky8eXSSwO0yP6J0x6x3gFUWJzaFuUe6RAluaRIFMRF6x5n2Hrsd5oaedQfEe6dJZgEok6jlw+
MPjN04IcVZhV0cYmRDfUdvWRDrmtpykpl5oNV887dlUslv5s+7s9A+cVFG2fWBzk3sA/piOtBkSF
ImxWFsQn0SRO2rJfWvDNOCQi81RtNuFMjC5Bjh41vkJN2qgDyOmx9QXDw0POx66+msXpEXPEej5m
rrFhy3KBkN2WnlMD2jbFd6Tqspx26axQldMXnnRd1wXEYM34EjaIHk50aLjR1go2yMPyJKL1Ysz7
8vW2WOrvr23FWikhK2Oll1xDt/urXYyc9tBexGRSEdvDnPg4zZOBecFh5HX85WySYPTAB/R7SS9l
v9oYupex3ZvqtWRqAanc83iHLFxmV4jqmIchg7fQ7miPxs38C37b1IKVZurehMtBKGCxtli5kET0
p/aAkn9N+Z5bCOeYJXcPP4IuzXuIQioaGmGgiu+j9IBQ1dgxm/E+O2YDjL5Gnng9P80mV6CihiSK
CUfm7v8PT+njgXb0hej+WaVXxVXRHfFiDkm4pQgTQLAoIzLV08KDfKP07c66xO9xM4O0XITv948U
M23t9skb8h8AOVfFq50A7v4UJuxB6mbHCuv3xlzfH+gxDJTBX+23xb7mKhsocFDDKRg0e/iVlgua
i2EPNbAhDc/ngdvqEXSzTiti6QsXW5B1a8b3Pz5TM+3VFvZV7iIFAntsWRXM5Oy+q1F0yqY10mk3
x1dHxqPVkgitUZo9mcHTLU4LseuiX8OaY9Dr8oBYAXQS3cs9LKoxg5BDvoUyeythHLKOQ1tteJBV
WT2tC7minc3xfQQQNKfD1rWmhoA/lEOFkehKe86paUrszS+tczUieSj9VER1wdX+gOm0oURUqOHz
fRgOKL+W4kvM0aU0h4n5socuM/vk5ubTjTAiBMYGfnbOLC3FmcQq6eSAPV7UkRmWcPT7LM4HjisZ
heueXoLHLiz1xDGYueSCp90Fx0JdccSS/b30zKkldhj+mJutqicr/tt6vue+VAoW7BaDSy4bi5xc
rJbZPFBSplV45gf5C4f2vdNzIukm6FPN/1PFR/A9Ibd754zcaTOeyfWOVcUwzcMg+InBdiPoEG72
yiiHQ29/wNUyv2zV1ASKT4NN/0ajrLyY72nVmyng4V0PvUI2H9r6PQ2Jiy3ixF+N/lQBmfsLRGXK
qlgNuZcQ20Iq0jBLokAlArN7DHi8KErOcowBb+R2JPQirql5tbzQlfiOSBd4kyVR+BDGgaB4Fb/k
rYw39PtX9D7UGm6eb3codc9gBp6DJJaoFvsS4n7hCrWvjic8cHrD3mrAH3uiGaszqwHLxXwB/eBn
Lu2dBTtfH9sSb0GiozNZWpz+1MAV/VELdZQhD6YjFswPhvgBTBJFh8/mW3VV6MhIquCwDdeXFx1G
ShsZizxTlYE8WJptmwKqa1tDFdJSc9JgpnXK7OKh7FH4YvUVT3V7XO5OWRnpxeuYaeaRT+dQm8wj
5xsquyRQn4kfPkFBfhl6akzPanhgInPJEz4VNXIsHWAulfTkzaRjvCmEBV0BrADAJwE4g1yBUYVO
KHAaMoKE23d1y6mRs2M2k2Ax4dmyvNHeQKGulSPEEcs0lwgkYpcW0CLfyey2nMrJw3XI7hFwOKs0
L6tzXJPWSn5TQOwoNJEwTxXWKAP9JS6fU6/NZu8Q76sC1VhoPgqSBraygL7+soFbo/b09/wf1qbo
QHD5NW5ShivEzKI7vgFfxyjYoLSltC3/qZxdV+7lkMy/ouczpbFT/9IG7mBTyNtuYlQt4xKA5kFp
6osZ+ipbCW+iBe2Fc4euw4E6Uars/hkfouepRHdNAeku6ph2Y0tqtk2dq1E/AsOWAeiZfNjFPQT+
APZuxYjdPUD7vZHX7tZ4pgA2dqfbDMO9vPCdFTd2U/NFnL4J/X6v89AqOHFn7V7JuA/8yygzxYP/
jJsSpwEZmVNdoleAxkX97Koqfnr3BG7oKwuHO+Kq/GDjkWL6O4kF31vS7g6m3Cq4k9XKCcP7c23U
ICrjbq6A8YiL9jFPk+SgSptM/Gd0eOoJCh9wCvQiNojMmHxuD72RPOleA0acwC2VvcjDgToPr1UG
Ju/0P5hWJY15cRIZrH3KTMG+29kGtQDwBfkoQQrcrLmSg0YzaFLuh2mBbd/UE9miwVnCXbDkzGIY
/0YEAaYHYnbxsQzAFHi9jBuP2n7oY6KVvBquGt+PLPl3lLnh0YHZQ7Yzu9Bsus9C3pDi7STCQcSD
/bWgcj/SUAj9gnDFSKiqN7UCykjGK0vWVKDZZb92fUo5T/5Q5eaaG0tPbU/EdnqZ5lVIbOSPOzIM
+Hr+nvOfRj22FXFCL/VFhiZZGjl5mmC2mjSRECEHIuVKv5N2wHYl5q8d7IcT7yj3THfRUI83qGea
e0gG1XDVxLj5cOuwr7VslGT2ZxhQwny1NMX9J5Qxa3ic22YC5U8maiEvlupu4yEbps/ZMht+lrqs
DDp3bYeVV4hH1FcBISOnyiyC7uc4ieBnHTKWLAJcgUE8TWb4UXo/OmDJiDC7pZ7J9zS4dMiIuUGi
cTVXwhjOocj6MRl4T+2Z+XBw5fHdv9oHg2yC4LPgOrKAye+gNeHXOXdzgkQSl3XqKmEcB6znzz+w
VPA/mZZdc8XLxKeKOm+HD+QUV3m8bcvqWzjjFlmeziCpNrSX00H82VfgKXvGuYQi5ZCrM+lpB58l
xZqCUdg8jVkWpcRrw1X+mGXHgnxAjkpuQAWAN5GUo6ym2gzWyUHq/4vOb6mYFN6JDnoSgagcwPR7
dZ7AR5F/ypsispSwc/YfltwWxz3CJ1V0hX9J7jI7NiKIxwUVyqmBue7V1rUfn8sh5KtsZVRoBFEx
Gxv77IumsvDjEYejRQNt6lC3x6zeJll8ZdJRLC3p8DANcPoXxcvaqcwnAB1AQQFvSX+G4udtsdZ7
gA2BRC63nvQCXr4Yc7khleIjN28yVGaIADO4Y4fGsiHPvs1wWu1AZArD5/UeAZsQ62HHiE/1yzVS
A2BddygFcw+EgfCeiNxaMpGQ89UsYoqCL04tRg9TF0VyUphuuzOx2xM0IlXzYvrdKnHIMpzofyAx
lF0WH9zA3NfMCb/jt0rR7hSw2lSZLCyQ14JusaGW59YyGuhuxuqz86yIlxsflfcxCqwQtcOBVZyT
EyajJkrmdR4OJuav12/MpQ45DTS58tU9fNBUuUR8q4jM6U9SVgra5xxcSwl5UzqpZxJPX+7y22dt
DzvVYQu+fqDcrYaLT/Y6aeqn2Y1Qx854+Cr5wKR3aJpk5Y1q4UKzqwy/4WEMc4wh83PhAUQlBPLg
SG4bxNEjUPkg9HZY7oz8uDA1YkDBE5ysF5UYiebKq2FHNAh9P0txHh/CYMgLphv+Zl5xhmhsh7x3
miMEEYAIxX44ZQkCa27vzbI2OEof4bVXuaICJHEmegDSpAik0BeBxEo/V9HC1He+TJXlkufdtI/8
qg1gMY3YnxcWtd6vHglpraSfKw33v1+Rzuwk0T6Y6oTiaYOCGfhaEnopBMUwikivbw+wkXVVQu6D
Y7YA8qGCGmbp8CzH+5Ixru33y3gw3RYWEGe7ME1ZNcqt1hNl3d3+uZ5hrykjGh4aiYwAH1rkyMPP
QOqAkDWGkaR/9IUuQs/7t91cxCFbiYWtN2v1ctpBz6OkwhdOl7W/us/yMYcuexjNYqKAGzSfnnqk
F76m0aBoTTj2L/QuteXj8wYJ6AzW871NzbfiwOuolmTS3tmJUJGDRvSecgjdS6dOgTbhTQ37Hoas
SqkqfVnzUTVjEW7mBk1KGs/iXy3eBrESyPWxTKFMM2UpvdtKO8k8ZpMzeG7uTpG7HqkLJCQ76xj1
NJgCP49PuwhxNaeXVmbxkUieiLowlcdcpJkAIX7ffKMsgGK3oJAUK5s7kyqUpCVLMOgOgsdpA1m7
yd+UAo4ohhfMMghdMMOkeNGdPhLVNvjgT9v8Xcen1vyXtNlHpWq7k1MthEsti4HihpqPiLus+2yx
zeKOqJ9E37EZFDu8KxbaqhCHefEdGB+KwiZtP3G66szUSYmqbEsg/5MKsT6rxXpXZXod4epnI6AI
jswgVIY/7OsiK4aWwp7WawM/30omQYA5APRGPIIJwjPLdCfvRy2nbmcCcKIB38hMpRig5yNlnMkf
CpqVHbWFLbqe9yXQlLBozQHW/m4W1Vx3jOx5t0Jhsieb1CmZCzvxX4yQtmAXuDFabvY7AP058G2i
zRvmmto0BUpDwkI5qIUDSFYfKv1rxjBDooVgjAF3dyJmA/CkNbaPhK+W0QPDVyxwTGefaWgH8Xqp
el8QrGVjNDQOyt24yHe60ygsXaHYlcDVreCXU2UPgWn/S6IXjyRNhhZ6+GC9ntIAIyD+A3g4frge
Fu/MfxlZ8IkXdi8yTLeFieet7bLTaPR9TggfubeYFomViRdvvAg45atUlDQYSqIGU+MpSl+VmXG+
PLIz8ymX+JmrDeMBSWDr4MmeV7bkbe5YFb0Ul4yDVnf5qWwSTxEOLVjAeYZVJD6DaJzXewzKJr3P
iXsExTLFXDxvK8ZRI6tAPx+kH4Wg3+WhK3lEYuUjN7tm/YiP2m2N7BspUUAJH9O6mOMlUTALpB7Z
aYYdbQuB/0myOR+FjpuSgXDEoIGs1EqArcyklUd82JqJjCu3wamyyuckcfXfmHXySfoGOZ1MIZzQ
Y8lywAqO6l5XExx/8MRxHgYoFVi+BwfTy6rIatOFr1O2s2g9k4qjZ7hy8dlClCjYBcXeL88zKhzD
rgJUfAy/AJoWfjqUw3sB3UgYltJrin3YHrV/t+SoXcaNzE1IsNqQ921kNjNB9JhXjCeo7nM8PDsF
as3U4biUJtU9EqbAmfyVQg49RoYw6hITRuFSSHUd4+RYp3i/lIjPT0adGE9b3hDenoRRypqzMVKS
KcOdz8l4pHMFZSEo0TPzCCCaintRC/F8K9Srd2Enr1BDv8rpghnv+Hfu0hsYKuw0tAwv+nF9DOQK
cd+AHXqUc2fwETa3gJ7Dh6gKMituYYC1JrM6/vYQe3RpylpQ1/69rzvZwHph3qQeZo4qQwR4cOkv
hNQX8YdfJJELAZEoOOlzqadrOSeYMExC7bxPDjLfPqChN7qhZgGTLWwheKUkLEETCKpowxmzos9V
AdddBcOVkwFFASmNhrd9ixeH6NLK+xqoswgThCU1j6B20PGEuWwA6h1i0n/4CjN8gXH1FDNWE8ve
zTSCj6iDKovzq/j9wIu9jXlO5b7B/fZBxOvJvpMjDuiGLnE2AxV3Y/sOeTBVSvuhlktU6afPa7qV
nEePYKqy/R7Lz4i+FrotbpZzRCUOEkl2OfIueVTdYj++F4l3OCJbR1ijRYKPbvsC8WrP0OUYdqKv
wlbBLf4rLz3RLUvq6PDWrKJVDApFOan6p8b6ba4eMfWLkzi5rOAsCH+MxdaMUlb3Rq9wipjEh4j7
UosDMN3v+sUSGd6/DIuchHsTOhlrMCbsaJmiO74W4ARJZZ1oq789/aLb9D/k+2LIrkcQ2ggweWXM
IWNA4wy0Ph0OBGCUP4Z58/KhO4zuiufwjYAHIAflbi6rtHD3+cB68dE4XcdZxaRkbsdJ+sHYx4D2
enbpI0Vz0HAYgjeC/TndY88eSKu8JaQHt9+TioBoImUIsehzcaeoWFavQMKZ+StuxpvJgBfICre1
coEShRstp75yi120JvQY3lqP0+CEVZy/3gEHBQiiSQZ/fYPoXr4zMOfSN5jDHt+FWRC7KAF6KvAU
A2t8waaUknLT46OTYbfsY47xRiaAyGdjWKd/oRSzw5VCvrAgXz1pHgzqy4zKJQ8IpDlYdgf56FXP
ILsw/weNUgM+1n/JGpOGa5L3/pAykn1FlPRNxAQ/9qTLZ2pM8FvvY2DjdpctegHRzqMuPmwA76xJ
2R4aILiPerDjqrHrrn8GK4AWAWU9nyE3taH00sHfHUcNtc5NOfcdYAfBDI3hr46eDhyDnghteG3Z
tWLpVspKGfS1CoiO8AQzX6zn4lC8ynHFSY2rR0i6STFynd4s9GSyzo74HJ9+0U32Ow80MXVFCLc1
hf6Vi8r4JdP3tsyvsJEWJ/TqnPLk7Aje+5FkQiO9N/z8dC0hhdvjlAbVw4mSnW3WB4wYUeX6Phij
Lq4xm3UhIKrfZw8Xlli5mcrj/Dl55wWmvqEnPb1XVe6tRGQq6hJAZ09k6dZjYA43oYcrylE3bR0z
iqJJ53B07CVBvQWUgm8mRBixVK5iphzvc9BWnjsnernZ9eFx/KoF6aGfJ/DKBhpGgbrfuiQVCJ1k
a8Ire8YbQ+sseKtw7V+zkZcMHlEHuLa4NJg+l/TnY1NWG1Zky6OZXISG46Zl5DDesoXrTB2mCjRd
/rwuHTxSObv3iHne0d17h2jN2gSQ4A4BlJ/PA+QkDSBICy/OJi+aardVkfLEA9dsm8Hj0c15o1c1
tTdb8ub4I4ZjeO45kKnWaBGt7CLn00CsOnEN4LlX21wErHffKpdz+LYeSNCmD6hkzi3yFAG/4eIg
2YRylKe7NQsuKUy2o6DAoez7/wP9OwmwinJND9bi3F5sGg1dZ9frXSCAKx+ObNAuMBXbVDNeupsL
HYk5M6gmtfM9Ko+NLjdmp1Mh2vb5bVE+gutBc1tfe+7AnkvAk5JCBNwcL92GNIla3m8EWUzrFWwC
x78rv6YAG+5gLb8McZZ0AoxfobKGAOPtmfyqdmce1aeR6OsZVH0gnWxEyDD6NJyy7Xbvlci4udby
E1htT1aWlvv282OEfQdB7itqymP4iLAHPrrcNFAXH1PW9WVrL5Pn823adUMUtHh9lDAePrD/p7ZH
WktEvhR3sF79FCtb6F8JHFQHYQLLmKPjb5Q0oMYM7ceQOc5WmR+vYsQmAIMehFCvVj9q6wNwGneE
lprRv51nVvfAa/NRR6V7+LCRX1UHFJG0n86wuFSCjZBpULYKIlznomXn7PDdf28taoTPAe3d6Ltv
B161gyNBHPq7UVvEKM36hNYcM4wExah1JjF+oSbXikBe8+RyizMTCW2UzuK+GIcHqZg40e3UkmIf
FkjAyt5D6N9GJJU++VXybQ1+gRfyZn1w+xg6ZwuGeToAuHx3irKgAtTustjs43k8vZDhpWSyqf5m
zK+weIuc3WrhloF85hgINhfx9im3Lf3KIddahlaUgvVY7tIru/CBCS8rhictbLrI3g3lGoM0rqN6
aT2QNHhfBHvXEgf8z5srSmslQgcMTQcwDr8sMuY8zrBm5FNqL/kKY9UyUVJRVM2O7WqLm5TLw2FV
il+uovhj06C0RGn9b964Mk/XQs1Eq94mvGVDRvqVprFwsU8+B0JwC7gAkgP1NV6EGqIuL0N3NI7R
fWC7H28Z8ecKZiZ8Pb2e3oHsgLmnETY/yIN6tdp3dPUt3zfmvn7uGGpNI/WFSupiEe/B6uTW5k+4
wHZiMHS1opwrzTb8NZOVWai0jVwQQ1HmFqWcVjxWSE0HVo8LlSCLLtQnyW4TNjFufaDWLuEyB15P
4rTFIbbeJRsLbkuSbMwamPQJr3aTvdka68D5Ep/7Zd2+zO/qCbF6ilUrHGzOuGO8Qmv5ko/AQaeq
/ivdq53k9r4x/0B4wkOwiOJ3D0EZ565F5UhrX3z2ZI+cOhC8McTlPmWsBJ/b59bDn6WECCrg5GEO
omZs/3mAVq0grcEAfKXiq1q6lh1XYzx/CDY/bQWhvtBnN5q/S344JU2nc6jMSBmcOMbp3HDy4+xy
Tj8cdtNwdlrcWeX800406gKWvBhrfIy2Uga/eEqhjfNnWqd9omQA/tsABQ0uffAgcINCbaZxur/A
Sf1tQiL/5fgErp7ZweEjjzdFeZI+dGcpHl2FCRuHWQYGqsLwEavPVeK7Y6y8F9G28k6QpuO/Kt0n
+DzgMjc2KMwo1Pa7STTD8uUTgvR8xCA0QQ45t7zSpG3CFGPVX3K7WPQrOkD399nueuoaj1k63/RA
eeBjrOen8+pfGK4aD0DQLy9oFHqrBC9dMZU2W4Yu+iZCVUdyCU0W/B65b9ITNq7CMwvhUB9+DCXg
u0YESO0RA6MPYlcEOt7ao7lDrtDNkhuHHJXoudBcm1sd14Of5Glz6aI63C9c53tFuWUWjDZpdySx
IfoEQiFx+b+X6WXidqjbi93ihsPurI1hIuwNzkEvavnIDagkObL5hNGCT5tXtBtrhlyaRjcu5vZj
T3r1vu4lXImL888aPhjF9U1Ejk22ayN+Kdon7t6S0wxUBBhdXPdWiXGfEhwron2+nDBzShVkPK0O
I5KbcWjx6v26dmyeylUrNiLjGJq2jaU7fudPL3wmvW7796pfMPIRFRD6hKCTHE4GiZICgtVnneEO
bdCluq8YPC2HWdx1uTfOXbiUR4RqWKR3b7scYsqMcFy+86P1cqUIgdWDSgiB0kIbGYv8ap4cTEj9
zs1pWCHLk2wItTAG5h9XTi81AqoLqGOAidZl22OkNx63j+YdzamjmS5imwkVh4epKrZB3D3PkFfo
pMLlpQGgCCStTnc+db4ow8LxjLhSQx/3aMSOKBPHhvmCiQVQR6FZeEg4OHIU3SdrvRHqg11D0J03
kno+6KnUO+5rlLiNxW+dLfvNGHwc7IgumnJFpYpnC+VmUw1FhA7ljNipmu2TVDCJbh8PT4vctbsu
Q00I5vW6vQvVPqjSorBIioBRwlXuiOG77J3jH19yF1kTNTXSaXiD6NxX5QV1iXRCU84VTDdNO8uF
UqT7jTxAZh2/B2T6mmYSAjoPMtfAAnqZT45Z/k+mqEjDGcKzdcA9YRpcbX6hA4EN/ZpybOsvdkZ1
4HK1CTgUxK/JxanpRINwtxe393tZoTbU05IY89Zc0rLhzk+5/yGAk/wUfYq8dTJio2631tJpZcrf
oVFmduwZV3bM8JY/y8EbTFADFRDWsZedqzYGCv7EVJvJCZn5e54u91yAEgbMm8sw0PGtPlHYPXba
wMv9hY7AhPXwYowAaIgkPIZGYPqvOzc2s2peGf44HR0G/nS63zoF6MCY4b+NQ+eajLLHUdd2EzFY
9gVERSK5P9KaZplG/31EF3+v0G45MgYx8+jWr/4D1TXDe5D9maF4eaqChwVEIC6AfzXqDSYuhPPR
5uVkq7oRliaBxddH8uzFjzHHeFU7RXZfUoanuFwRuN561fgfXtnfm1LrSUn7h0t3TdNETMd+oW0S
uxlWk2YoGy6eDw2PwT4alpw78Cb7c4AsYmcgZYWulyFlESeMh2iZNFiXn5sKHRMw3DzY0LK16lIY
lJhY1y/EudhM+bbuS12e5aIfJOgxt4JBstJamIIChYvgrRnmapQd+YmtuFOL2YsMm52y10yIAp4J
sEE9OZVgrBUKEDWIekzQtwTzPjgMk9gvDxUVJs2+Q+zsPFBDXLF+f9r48V33B9wJ+gdQZzZkAV4h
bh9DK5tmnKNEVUv5V/9Vci769JlFs4NWClD0QZm4Ccoo7TWhJNZ+UqV67WduGyJzwRHgf97GL76C
H8UHWecAubUeC0pbpvIDNoKeSkOeRCnCmM/dc7IVNg4XhFWPYMLvSE1r2+ZgLrmz/9D+v96FZPUd
DS8Cn/4STmV3n4WUh558mmqRY7kTuXwWH+/VMNEYP1gHvmbLuk+EBTFvzBaBIbAzceRNCYHfoTzl
QQ7/Y5d4aexdzpVPnEEZ+bnC8EuFd4Cv76/yMNTuNCgSd2vQCvLtb13yvqqhr4apxXrB+mBIcIae
1+I0rF1milIlTukppfVeLDQLrcptqRZ7t5aENX/Syo1ii5iGA+yrashtscmiYmtZ97ukMUZpuzQs
A388V5qZwnbDbA/Unb3cdh/Cx2AuRxW/cMEokAjhH0tlRAPocJKsz5fdRZH+RkTj60crac3Ko6AW
9VOkus1cD9DAruA22npO30+RBXW84Iuos0lgsVb0yoqSeYKoMdLbW9fiY+2dfILb93D/yYDZTLza
WD7iSqbOJ0vsyuAiqQfAxenMd3LFF24mw0V8GqzxK/DbJ3RIcslJ5SYzTYPe0vg7hEpA3LE8fWRY
Zdf8mXhX1AYefOthkSLoz0O2w2MdjakJyw0Ipvasp0ASv2SzBTPKTP6doUe/lnsyryapHF8Ehl+U
NMvUWMkWiDWKT1Rp7EJ1jE67BgEK0eoKHkvt9mxTTgaxvVy7aIzsPM9VBkJec4cGrQ9yW+qElIb/
4g8ul6HophmMTC1J1UELEx5jX2Rct9Xe/yKJBuCevVLzsEfBmODWZ9MfXfJV+GujzZHRfqKvRgmv
tsLEIfKjczG+YyLgJJxYQlKMABmEFB1YJxy3ndF7T00LGYyHrcOJoNXXYtkCBAF27WSztjw/geb0
uAk2uNBbXjOXymW6yodQKD+mp63Oy0FQRm9UfjjhIFaKQtb60IXKK5JisYJ8bK1Yc6vB7HiDNAFf
qQkLU+E/SFdCWkk3S9tGnDZeRMRfAz/+Kf4AQX0DghGYU1j6Luai9JqOXvGaBbH1G+jow/5AqpvP
8t36OgAj4zzJG/yppsIsT29g3h/NxDuMEfH8bZZqsWCVUUJyZr+rIbcLwxCtdXR4CfLSs/xLPXTG
UPxAb6K+IaRl37XCQe9LS3+GyVImVysPcfUqki33TL1t+cNswBpoAb+DdENupAZ4BhBgA5Vufz1R
6ksd6CgQxjkESLGdq78Sw8vGbRrpxwB2gMVtMO4uz7D7nQJAWjXaC5L25XDfGj5PlbMAX35A46xz
lSDnJ7Wa+anv3W9LBjollem5iIKnTofXAQ+VUVAFGRxCBvTITkRbnm9xO2Uv75IA/ye1X/uygn8x
86gcABfhIFO9R1Tb3LNdriKm/QA1KiBorVZxcs/oRlXAbgsSDO9JRkwbAjqZnymqQNnjlZaeEo1u
Jk8kMBmfa72HonxWRDxL9zE7vm09Oqp75dqluG/w8N/mLwYc0xTX2bItWfR+Jl87mOPcbJUtD2Vq
zKqmPy116OZOLLI8Ci7Q1ezeI+LN/e0ZZahc1BoXvpJk+LglehCPAg7vS2uetnPSA2HIlz/U0Qta
Ew5tyLFxhvLJxA0Bk/rdZRpJiM1YG2GeSc9HmKyFFhBLdRVX+9di1+CjT/IDq5R4ROvDConWSBq7
gADocqji3a6Pz/6wQg9bBpN5bb2W0WPseslupWpcHCQrKeG9yjttETVr89nl0Kkr4Kyuw+XO0zBG
Cr9grQ/BFhFJ6GVtv+JpYU0EhmUKP3PjIltfiNtQKz0mq3qcqqt2tgIn5m3lRRCg/jTt++Ml3w6Q
yt1c1gVQeCpRYQzlhn6LPX9IGK+WkdYCEPRFE5pPL0lSYN2Yw2Any+xegJgW5RCR3BIUY4cddczH
p/ITxv/gfQujAzGAYn3439M3PT7wGPjGJ0gtU04cLoYQc68Jhr8IFzq2Wx51nq38D6qZ+x+1Piec
OcjH0xxJXVi8V+FlcceWkFdPmokdRMm889UtMvk5wNsD226seeZJKm1k8iNF20Yyxx1CYz8/nzls
kMwc8ahll1poW81o8ULTSkLph2/BW03kKX5EK0d0jkJdQJN2Xo0fqJf5I9vbTKvHV8nCJ+7Bs4ES
1br0UUDDAedzr8byvfJbndrLmZtw3quO+V/P+6gGHWcNZ05S5i04J373XcpXxuek0B9AauIC3CE/
7INQvVLccwBhd3ZWDp8JLq2tdTVOatcp1bIPx+JdupoQ3Q1vNrMdvgAlBkx7VNZMX0sgI2O8/isg
RCuPEZQtD46zKQjJod+SX+4E13hm2SIqKBjFNe5s0icwWCeU+jTCuCLSL2mRKtJfjKuYSxwdRNmk
rl/YPvMsPBnNPb5n5AZFJZFOd3DuugYxv3IFyw4i290k3HBN1Wq6yijdRekk7jjssCimrxmO2Hvt
Hn8JglW91ydTmMVBgiSEpdYDA+8f+ljl86w2k4UFHiWPhC5EunxWnvPcu+ouytOWZmq3EL2kb2hY
T5pJLWCz8OecqqNX/hy6+8jLvayhdLWQ7WU6KUiMW2nKau45lKtNAcKPHP9qFVwKTbW+VA9/1rZf
FBA2/kPbFT15kCe69ZrPu0o2bykZegmljlqm8m3AkYiEfSMDo7Kn+r1GZFobJ6BHfkQNoctfDnLU
hIYq0mIYGWhnBupx/GNRAPzo6tMuG9zV65YcUMe8EkGWnuDCQvMCQKGvkZyqyH161d6sBH1fgXO7
QSKd9fpplOlcKp0Hjm0CD7giQE72FVxy0ycA4HMKNz9ybGs0BSEHOa2wjXQrd1eW/ZjT+Pi/qHdw
NvLLMx2ibj5/0wpdknyq2vEQfuY9KqB350YpKrJJIUcPt9ZTE/aKC12FQ/8a47pyUWvRCXu3CL4B
BVrI/1/y9XG4p26Qtck5EQKVjzKIsKcCzOWhJynZ2tdcC2vU5NxnPM+pB+q08dcyRcJNbTfCgoL+
W/oOcRACDJZuLvvkRTSapkuRKvv5mOR4ilWkqJCT2obqBEKUpuZfLQtArtV+5SLcy5ue9fY+H9yF
SXAGIRh77uTHecZLrc2fZaOUWxI+qC7+IOSG7/Lv7IIlCqUNLzim0W9KtF8Ye79J6NXtYgdZMI9E
1HSpDPBHm7+zOOHm8VNNFIPZT0PYJYLjTm65iynyxkkoYMyS6N737D3UvagWT465O6zc6Dj3/Cct
yKFHJ1Jl/WAcA7l1ehAOf48ZMQIyLigkI+0LZEIy/oGD88v8l2SJpXhQmEd1FBqrNidk1Lvp/Viu
5qb33Sd94V5Tk5kC8SPnRlBU+UiKnm6sBNF5CdWrGIhsY2rBDPnSydnJeQLe8GUOUpjZ3ITNEYCZ
nsR/cmrfLSkB3J+uNDhaIe3Ini7LEpf67BwrzgNRODQcYLxNEpxUNGvUo5FNRKGnpq8RN18rkNDZ
HgZjpLHMZIvRp9jEy6hQF+jyhKI06CWT3uAsBl6OxY2L9x24yGTKg2A5uYx6k0cgCgzldA55j83a
sHnoBbb05b7sE6CzvBrS+keLKH2Mph/u5/tFt5cBj1YqB40YJBRZi/cCWzJ5A5aLK/Xubvxo8YCE
6ySd3JyZZ1aJNJ11gEffTZZOiuSddmYIhHgK4GvunKB22b882f48GjKOsLBMalE2zY/KEIZ48w+m
TVn7DUeAfp794FzOWKuJGnIsQwlgeNHLeeX0/8JcEDVzsJC8BDGy8VJZ/PGO5TKfFVOSU43sqTvv
b1mz8WLsqhpwWFuuKt14/zAqBNfIVEoovU7+CZaH0kq/sgh7nNht2dGGKk3J7S+RMKnG5EVkSq5R
e/HZXixU+a+zvO8fFEMxJstiPEk6JL0f2NfDccHT3xpnzid/Oklr9BTvQXpBSiMJGYwQQi/JFSsi
MUjMbeAWwGTdvKdOxgRajb6hMJFVu+bUAtT0aQoD3PAfoQFRGnVg5kZdHpAWM7qZqPvvKQcXnQWK
McUdzZ6gRjhOVWHnCfF2WO7WlUcYcxv1n0JW4e1aOlRQNKqvac29z12LjSgueedR/e/+C69OwNzP
AQWetjw7GaAqpL6tE73kS03fL2nRreHXosvwUAOmugEGUMIzOEE5orMuTdY8L9LszBSVN1Lss7sm
HoWuGrl028bSt5gBP2366Z7Ph8Vkic9x1kR6+FVtxfa8Z0hOwpFQStyoYgaDUIl2lkshSoNsNpt0
WbQLWEy0esacwr+Ut27FjfTHBU6l8vwLK6u+OcnSTYhq4ebMEndxVgn63nHxxcNPnFU2uF9sXR8i
Obcwk6bdBOi+50KnihRFpbyKR3iduD7YGJzBqOH9kmoUGLkPWN3BhJM5bA+n0c3+VhBLLFcq+bNC
CaNrDIzwaxrW04Tg0ayohLksdYUewKQ1J6Q9luIcM4u75DsGg33e8oPLHNbGqmkrlZbsPK80ApdE
gyJ7TSgbs/K31N5GoCLz+d4mNR5CFfoSAlwHU4OFlNAskQwQmBbCiB1p0XL8iHQdnsGaAN2E2Wsf
XApUul/TS+kYoHE5PnE6YzPvbHRxwSc9pvgwj2RJSq0SSvmh//Xh4IrvsVnoU6i9GXka6BskFPJ3
/lelb/Q6IIvNzkd/IJeoqOr6YJE17S5vH7gfK+56m7rBEr/d8mzHX8WbsaqN2lMB0SDi7YnDMo6J
aFRU0CGwcddISIl9wxovkfxnm38oTCPy78Evk2DSIE9Ht7l4fNUlccNsSiCX9s+dB3pSqxsifRR/
RWoCNC8lH0C0wPCoJQC4YM0LrobFpQo5aMkKKxHm0xiRPZJZFCt8YVAfSu5IvOcuXu5tIy50Nr6Q
J3ZYUkVXmqTHpguE3itvPfcnK7OsUWwLfG/YxHH4of1EPtXDi7c9tBInNJ26R/PHPl4AxTRD1u8e
BbzThwzEuK9Bc7t6i4GS2nRJvXLBUlkRgYp2Rm7LgW0W0FlcgTwAGxCg/RyZjlXKRclMKHwsnmGO
ekx3KbRQn2c3AfLxo1belpeOTWxjvra3S5aENEMXfOvfkoZEi7YYzGRVCsHlRWvsa9p7o4dOEbZM
VXnS7bXZItMxh+9P0iDaO4DmKxxbG68g2wdU8qJ78Ldd08YA86RToDPfc16zu1Oh/oY8EGyKkGs6
Zh5YWszwevXDbtqfnkkskSj83a1DFRVsO4QcqE6FlEYYKJmNJ+866c66/vD0HdThvVH+kWRxVCpL
1rD6CB7EoAuAa/AKwX7K0aDKwhAIZJ3cvriN9kznlq7iO8VWZvPsLlYa4ZemgCRwIloCTRth9D+F
ecqMlroOsWrAhyWFGCyZmY/+kEZAlhJ16DaHffgLzj5DorzvZX4pdxGKj5MKTn8nTWluhPBs0w24
sBgK7ZnbtfqCjSOzoXgkpdqiRIamA1yd2tIbJHyHrLKcUsIQJBo2olDI4BMKPjcQCOpVflE/SdzC
S+Kt8mXWpBgBWpUYOvV5QBp+R4uMAxURpJTNBB1bC04qPfHB4nr1e/FVgrg4ORggFRfA9Vb6aC9O
LD/lrdqlOcycCix2kgcI3GpJ2qq1ekrt78WOhV9BLD2xCvTDgCg6X70CY9o/ze0vKuZjjWunIwto
tzATIe8OoePnPGoHuorAEIy6cGdjYF/az/wFLdF4os8/qa6RbDdGbGlLDmhyGA/pUUYjB0EV+6Dl
QMRPzqu//5VE86B/dmMpp+/sQcCkXOEu8tKlSYbmRnWxGK+7VIVHtjt3pT7/NiyXi7dICUVHJpC1
TKWtvnGG/8dNXJA7eX+VkssAF2B7idkKe5nXqNPjoibM0xtXWMHWKth3D6hwSeRToq5tyNMOZsQK
jEn82bxGu0dRVWWlEpWuXJmG50eIhO6OREomQVWV/gZ6CgUksyfz+823zVOl07B0CsjozXRKwgdw
F5ch8xeJEpVuq7R0fSaBXEz0J0pj1tHyPPSYsjUGVfS+Mgo6mZn1Wwmji1GH4VzS2uLRRzGyo8NE
dLqQ67g0Imzo8K2iG8TmV9PZeqQ2Aa+4Spbv0jOJy2BN7x38xVgr0zup0S1JOE+OEXazZeO9G3lN
+4ix8UTKdcuuM9P28iSl1Tq8RBWIL7hM+h5NhgQDV7zRy8XqerDugbvecfcjrngFgeLsdzHJ/Pdy
f1U09UgRj5gtkRDdbbTWZpHIm6vvaKdC4Y5TujajsD91VPYuCi0F0C8cgcQ6vBeBy2LiL37X+8Rq
XSDTWIgJ0i6KAz4z6ljHtJ3IdfZ0swuWbNP03qPpteGZvY0HQXhP1HZq2lRdK9W4o3uhIS3PY7GB
9MM7hC6WHzrnNqvUgEvz7BhUKjNsFMzph87dUA8aC4z74aq1uRDQkgwR1+8rUUze9Nx5Qeo5Jk0m
rqpJ2Gmyy1aZ0sN6+zhwwi2UkU3Kv1BT1oEs2Ae6G/B3huZaTcjlfjT/AYNNKrtqUxDbMGMRPoR5
MeEx9Cf7ZWAdSJhEi1Sac/4aKlDNYgR94of45oWgSIrKjpiq+CuwbwbNtZkYPhpVBIKHQKBvwchA
i62SF7ntuxk9dCSuuCTLaGI2fSdoKqy5pmt9xxRRibwRGnOL1WI5AT7cB4XRSwZYlWzoXS7rzYtr
JJB7STySGZwMyAq4xiBm6+X2nAIRm5gfDbqdCFHlfr+AM2k/1CVzSRqGbtidu+JnkpkMPZpKj7zc
eG1fbqRqqIiRj2YsMPpy7U/TSE0tXNO6EcS+ZppWT2muDmZamxhpDYAM9EeLz+hePVzGhvPJDng0
QzldbI2KGs5janwZVSB9mOdr27oMU4j1cB5B0dSWatrbmGmYqUuyRRGUDBcFLeZYHQTEzPyTkobZ
EcIur58Md4iYiEhldZs7ai4K2sYnmQWGuvIcHar3ThVQBJ6SSsjW7vaNdU+/8KYCdUZw+OAgJ3uu
IupGz65hPIUNsNmuExRvHyxkSw/chOaMX+avfZne7k/LCTSKBY1y8MHRt7CaqwZvPWJciuUIOIuS
mj4Bdu0njf6j4OWYO64xn68Pqfb62m3M8X7Cusnvu78Cx6b/grAlze+cWu3C3qPtRS3HgJp3PUc/
sN6Gl1EpvtC4NE4ah9pSI31s0wz3rvNQK49EaLh4EnqYHQ5fTz47xHpxn5aAqgpjT7uhBjiKM4sW
JyDalJ3s4fFtlfFkE9ud5AxTM60SjGYt85I5Q8kUbyqw7h1R9b4rXjr3cQ/Kyb87SwskYINIddJB
Q6l4ugoFLrZFZMStAG3U0RRflPHFlygRKEYSaH6+cb8SuF+6TB9XimfMezHbMIWtPKJs6JbG1cUc
wccWAbKe6TBOc1W6W4/zAnTrehxlX1MYa0n0EL/Sf7vz4vPUXXT2su9TSsBwZEywCw44jRuuFsRI
BwLCi4gRi4PfJW2W0Kxff0wOFRvZ5eeKZj2ysh5l3gwetJP3XOoUMy3qc0MI6/Uc481ytOnRwVwT
Lyu0jJjhqvNTxftPoCpC/SUoNsRxYSlOJbCdHAM30nCbZxxn3F8iZOetlI3YuoI7x/lDCEk5sDnC
D54XKZwr6jh/CMFe8Tnx9u90jqilXkX5JmjlsFw5l72iJPpAFjKk5/MB3tkRZKeeA06RofNytSsq
7OEqOGK6DqGjg1MCyJlWY6cNJrfqw6i7qa/ArHfGppLti29oM+m4/+AYikV8yzX78lzMyy4m6sgY
aQsAtS/ANdl34Ju77SCjJE0yNKASJycplQ0iJgxKOzGZt9xGkDIJ0tpKgDAg/FZXInwUWGqX54IN
WJoyXyInOGxjcRz8DqQd6wtaPD+k6JL+3gzuZhANcwCjn8xnPm0vRmzb7NHVUHLK8wpZ94ARd1hz
tsEi23SjmQ0/4vvRzItHHqYsUG5dC22rf7UjGXO9O4acl00m9J+2+GtewA7ozTgybUJEQZ7RRlpx
ycIJt/5ZA/a6HcAqixlREig6qBOmmPuiXM6+nwsv4PuGHW3aXIkI7giMpbzJMuRUhsZ5ZCPdZ/tP
wsoIKASTHGRlzNOBu/XuPqgz7IjybRlSUDWjZNEwjSQaDiz8SxLygvzIHdtu0p4o/nPMsWt2l6OA
O3CMGr9MAdMtxZvp+AAg9BxjQMoOf/KQ5cARzLY/+lC0JldEzeSOs6YZo1TbeKqKcjsDnMO/BFSw
lnevTu6ilzYR2HE02kQaj5/T8gT6FHlje/xcTaGw/mnPJDmGIdAToJ3w3evJJMkXZC1wrKNGIASq
FovET/NOXr5tHffTvlSs456lkpquCArDTkwm2tf8z07OerAEkyQOiq9JY7zrVUCuNG/NpFDsUnQ1
cNoHA/hSAGMC7WHwUt2R9hE7FeX+NrQ28pdhOqtLaIwsToHh7sKO/oBNLZxag5LAz/cv17xh1byq
g1QU2Gg8EG/JHWYu1Ooy6VdVEiR+eUO1+yeRPOeyyXSRDp/T+ijWlrQTL/7oHKE9O3zpnEYsh0Ry
rtVqEy4Y/U4CCLiherQZMdx6WIgDt8Eg0emw9Xo4XiWeCkXNmgBWgS//YTu6qAa7CaSf/E0uKttT
rz8vXoAXcTyLnGfV1qOKT3FQX3J2RtzhaSRHJ+g4oicW47EP4jGFzDVY01zWf7aNJtS1HmNbrZk/
Ovg+NuiLv94Ns37eU9V9/NI69qm8RnzISVkeCATUsNOr3LI8IIqbTeIAvYqe1DnyfSvGy64uZ17u
AetXuqs7buMR4cMZLfpv4tHAzmp3NXXHJ7bzEGrD3UcASibGU6SWKBEeX23QfwjuZDtjeYq1DTTW
0XCuAQ8MBnjQ3r3jsIY5bWnnFvA4/abaJLEaVI+4z8IaOFoIJyiGNvbwNtm0dOV7Sbupk57LQlT1
u/PeEJlv9mX2IjQ1qQ5eKi1NK3bKQxXT6z/8FDgDGwTkEKipkr0TFjKzqoc6VRPIanXLyb6Zn20T
jgBy/5BRBX32nFbl30mPJMqbD1wH4lx9vbYHjPmStMXyEHVOvhnuA7xrNNdkaIOabs+w6qa+9Cgb
zMwIAAkSNtBmilqFvlzoq3zoxIV9ifE4iFJh6SGnfmTVHVYsA540slBH5ObBBwK1SkUGFGpCdAHN
56HiC33u6nTjQo3kJQTSUEeyvgoAB/P3Nr4LCcVg9/3F5gbtKVLHvXU3to/Fs5jgNi6rPCtRTJ1q
JlWH7DByp+cTQM77DQY50ACe65LAq/0pSrw9J/0niAoZ1zqQpHe6yjhlewVMXSugwT6M5nvv/jZ0
gmgBW1UtcQOnY6A7Jz94bCWq3BSXlSeGyUM4QzKiQX+DQs8iCOyG46b+X+KZuKziR+P7ZICKgIA3
WLQpyWNZTt0eG0zUkYj81Iy6M0cfLEN/wyy7VBF2WHnIDejiM5ubkLULhJZ5a3VzQNjko7XUppa6
aUfZbGj6A4MY39SZ4+CkSzxXfrSrYLmCzElBqO/0XFbYaD9ZQI+ZQg6n0j4SLJJxSR0nCIFWkcM6
N8c1RoGKoxbn7tXlrExqC/B2Fd9/qGl8l6+f/X3/yKlTj62OWvSl7ks2NkRKW3ei5BFRkhGx1eqv
ihfst9cPrURXBDPilQVuFSDXYeByhPHB4NAFP9y3AiDS08Q1ot04dAlKWuSNwxYwa0ZPEeLz9hzE
6dK3orDJw3BYWzsZOZM6+jwmEJ4g2PPEGMN3b658GFQnoZCzSziR7CZyZLSEy8YbHNC3MvJjmjzw
D+JRJRMPHfZkitwr2PJUvNlBuuIkRvTUCwTxuoqW4dyhMIwYu+F3SUrvh/Yq0UqbYZea0e56OxbN
U/86YwD4zwzMr9LfnhYaiL1AvYaLMuE0ZGoRmTcF2Wv2IZKZwzGe8o2ryvFPp8++73PbNJYTARvv
+696P4Mt2nAX0xjVAbbDdqpPR+xf17O+EpntRNNG2xUUL3hwwfyJxjL1U6bvDU4HB2IcSC8WGifB
VmWjuHelxF6DNWhZX/j5IKCphXFggZTREWsIUe2tbUeLQcjDWaNhLCt3Xt6Dkc2IQhIWlfr34Y9B
60TTVXQgH7uMKTkG5obmEUH9CHoUi5HaevSwx8y3DEuGYbY4MAyQIkFGV3luVemB3Mqn5pWKvMfM
0IUbOzgjL70VkiTmwD585YJKTyh4Xbwvj25SA5KiU6HmUYXxvuDR474RA2l/uVhEoaQwyZt4bpyH
Sn4I4iMzCNm7LoVg1phUymmPkdTXjImSEnp95Zi7Zl0WizAObRWtjXjYhJOmLCDySOt4oRCqsvZQ
YiwBzePCZgYjcJqTKf8Z+p02vXR3/MPGnySSUlSaLtQS7Wl0ml4fPY6vZfJ4cxeW071M3rgsQlfa
kVTAMyuVwqdrQuSKfFyC4GfEjaTObYg4jEFKoIrAL2S5r+/cNvCi85XrG8ozkGmMe1MU6+oqaWXv
L7Z7P4oiow8pU/GZkTbkkoX1PzAPt3/VLZDdQ9IoylW7y3hHyGSpNVqkNnfji4hQXNG8qtbgaAhl
sJlGjF1pG3O1VhEmj6POXCZpdL9izG6JThXFs9vZ2+apm3wLo6n4bXernBt5MDBFB5fonABeysGr
FQy3B5w7FEHms2/uN7TXFvwIxm6/7ifdgZ/4ny0x1H5QwGaDNIzefffUaXXWk2LGQU+/SyZNG76I
x6bJ/2ivQgLipoycN4/BqRvsu+sH/ODbdmLtK5yjwLWsICTi4uIh5pFLxT33ZVndqHS0Mt6fJJQS
t9vZVzV3Tl7YU/zF8wB/Zw7aveRVOqEwIX5BkUdz+gYLviNjK8X08XXcZRCYqp1WiqTQWwjKos94
kWJguo7ORzwuJithKkevNkpjdHEt0ELhV8S/4P2RtKKPTgCAhGWcDZOHFm3DkJ9H086Xp7KzddGY
As8mRw/Od0EWQBHn449xHZRnqKJJFo53YfBDuaWf2c3hGf/LKljd1e27IvhC/kE82QbLsr7/X88c
pSTttkakQzEbjfx6t+VhuQrMCefKnQXOrS3iHcqJ8J0pQOnANufc9u44LmlOxRS0Vd+cs8dVHrUw
iw5dN+mt4GM6jdXeEbVy3vNUsNAU4hy/85dFl0Swe8m1zY2/cNIJAtE4kPJ7yqjTW8PP/rKSoQS+
+njiuOQR09y/QLK344IApfxrlU4VCJIcFT9CeDipyA4t2KUITtFbbDS/cd9uYwKeY/W3s7jiZ0BU
BP2Cvh4RcqO584JJYZlhXWCpAnAxvyP7C33g9PMDAbDZ4pyAAfDqOfN0LrKhfYXJwnbO+iE9mHKC
gyP+yXD42vzb9JK/LZMdV/eWwT1i7A9sxcMpURYZf1lcs0zB70L+bbgDj6cX0PhABdLafn9XNUaG
w5yRpdcEbWjvxIx38EYUsXuEppDWN7cXEIsFP67PdAsBIbfLgdfyzXQmnkAreqNJTSpRecSAYPqz
rkmZDLA0Wm4nsXFf38ndJ9UowmBnmGFOKcNGe98TPLDlrMnYxtIPxpYs/teWn9bazvlX7aldW1C/
jSoC0u1QXP++f9MplcnDnoQSbRs68PuuyhPq7TRTsLBxYGGF37YJlZECfEYoKJahXQo+zKoMp4iT
3a90RH+A6KeZr4FXH7N7JQxckHyGgdcTMYt7h2pqyL25wWz3PaIkVl/kn13M/f4cfs8zcDCxEhMw
YN/9q2kG+MUK0i6714VJnEfmBnMhkAC/2A5f/1LxN+oydAMypIZRukUCqP1I2jMtR1G9vKC6pbJi
d+DIFM59Ze72HNKDUxdqP79YgvCfIvxc+A2FycodZsOmYd7mthisewzoYGzfIAeHRYGBUoAB/Zy3
7r4XnbH3bykId7LIyto/tcB5jRcWwM5EOKoItxTnOvoA6pKRENAjcVEGcQ/iXMxy8M7n5s0DDrRH
PRtNG9XnrfUafFn2RUsQZrj7/6Ub3Ylxn6lv68RhHNA9CElHtIrtD0iQlT+G77Gl9SGn7XwXlruG
Z6S7QZbeRnBw7BfTUT9Oial0gC30ojR5GprknkcJbWt3o+X3V+GP9sArGPHvOqVRpt7BXasLaYBD
JulcKbCpM/o/BFBM4hqiDk+9itjJf7X6wZmaKOPXM7e77iQRHVkMJ5+oC8zQxN1ocT1FQ5a2MD3O
fUIYLs8HLSX2z3OwN39UmF3ZhYB4t5VDGO6KUjV6HOCk84WZDutvCW2XDHRphEuIFIR7HTm2xgpi
QDlkxDI2er63/i8eVEfX71mXCYmYByk64wHUz7MN8iPn3hzki2KGYpvMpN3Uuhd3wWym5B+t4TjU
gvo9HWrjWz1q53UL77EfkKqdqvLHS18/u9yXXWayYJuDCdVmuG4NAVoh0ImUE8zd4OExfAETqt66
Zbm14cPCaKF6SY58IjAjpKbWblnpW+Rv8QCjn0O58vbXt8L06uPaHucML89NpTQuqhrb46re4ZpN
Z49zPCDZsmFCnq8F9nr7pojxwUFew07AkGn0hVkftw+Fv9NgUW+zP5bjVlMBkSOGmYnEhEMXcyyx
fF333q34cxBrcy+HzL9OIAGufKKktDJEpB+UDmAsOAC0R+Z3hBc1C9L/8+vEKfIwJJDAZ8LkOnRG
8xbjsFHmmSxYCPnFa2hqDKjS2SKsH4jBeoi/JWJ8R2YIqxpGmMBp9Vw7e9JMPjjbaub2j5qleLs1
3BqOodUbSaZKHTY0JbYodO4t1n3/YxDhO37JZOjGNLiRdyHhmilTe+JMUI28OGPvIgDviGv/A+Ua
OL9nNqJkPGxLqiFsbj+L7SxnYMjyWcWuVdAFVXLM7N8ohJMnGe2KvX2PXaDvIeee7VIcd0qp8aYm
+ZoVi9nCOjOvFpYsabsbiAcM7FjcNB7pCpiQV1hXv/ZyVCJR4zfAy2ZKJsBUlCGDn/DdPwxXhOTw
GDd0zXKYtLj9B7E+lUbyFsgwi1dERpiLK6NSGAkV3jkFeD3u64lN3RCkEatsAg4mf6FgRoBeNW82
+l6LQH43/38tLi2eWSqT+WeExrkSDvCIDq+ixvWw1+da8Oxd62zbL6aqo8O+3WIr13DSfwDlPDdc
HBXgkRYINtj0XvKYyy/gK2P0U0fK8p7NQPeTt7Eim7sVHOK4s7EpDxVdUzW+oIeZ0lHLjvz0uDyW
kdIUvqKK/bRP8tDJDT4031qACkTmCxFNji3DBxK+BeD+joIMVuR09JMPCNB9fsmA5/nkbiuZ2qH6
g4HYHUnc9rQSHHsGnq4b1HxQLqNmVahEn7RRSs1Mo6KFXp6i5wwyG0hZj/XLyn+pNyGN2Tvaei7Q
0g8RQrJLbyIxIUuzDdEq5L+jCzBvzMxEzpjVYIfwS/CwlTp0bbthoXDePr06f1ZqNm4+PctoUPuK
EsbgxpSiYJsEYuK5jl2835CUoGGUjIRg7V697tU+/IcT5eH0iLxw6RDU4YhHjWpxg5vxIAW7IR2X
OZ4IzUymsNlhxmVf36+Di+YWlmWxvCEnMoIaDPn+FZK7+hhmPjzTxVBCOJogBrkX8VhcgQeGZB+x
ABbPOPpCJvxQO5a9pa+bGRmm5dbYJI6lfEgZaVJ2DaF6f+mfFte674slmkZ4Icbg/4ZECwJsJlZA
f3bUTOAoWBbutBoydaZcyubRohKHP5o+rqXCrxyb1nu5o3jAWZUSw2QTYD6AfJL/4QfBnyOFyLuK
zuP3zhioEvMU01d0IUHpIZ4BpHbxGvt94BIVfbM2ZBQUut1JU9GEiDmONX9dxr4CCXw2btCEn82W
9QcOwwXR4swkyDEFmKfCKIzk2aiCx6vDjm9yMUIhc4G6dVpWyh/Oo18dTeaGMLV/+tYHle235iZk
OEk5aqAMJ5uBc+bhTz0nXlI6tmRluQ9hBcm3LSggKF9mKf70tbczIZWk5D4z/V4rYRaOQ9CSfycX
XJ+ij/uZuxyJqLT2Km6GlJL4PezoxvMiVTwwsgpfCXJgSNATRGISStDaK+Zet3fRf+eaz/cHxQ+s
zYCDGZ28+PA4LLoiRZkOeYUHhmFiPo3jZ2FWN21SzLE5/c/OQTfWCkF0YebZjCvTkaNKO7kf09Zj
XuOO6yAKxDOP6R5UvW+aHv77aSa1OvrbUOQGeJRXpudyS6MvZ8/d+I51TMV5LEtJAECUGD4S/LpL
K3L1r3E6rmuVR6nl8meXVxjNPiEAkk4hj+j8soUWaFOMWhvivM7PqDG0xqSPKJSoALYFYlmuWR1S
N8TTE/r/uAdtTPA+46oE/07pWBgQux/YfQZmynkmNFY4ricJnijMN1oykHFw+IH8HJ45sEPxwNZr
6+lHezWlSWuX4xM7WretS9Wq5j1HQ+OuFbUGI8ft/dTEMIWw0tLAqiZJKqWJMSoBTA6F3nqurWUy
iAAZY7imtGiskU+4Q5Gqoz7U3p1aHssz69L9SfsKy9MOiB0Nax+YmdV3Fp9cOGsWUDA+AYZ3jZMW
OgqI3fvfWiqKUieVO33yTBuy8Al+if5CuOy0bUzpB5OFqOT7PXM0JE5jfk8C4c+TLx/4qsltCtJu
CZnyJmdNyDyEyhWddjPK5AURKaO+jrTcMG6571smb94bTWXaJBKTKq86DLCqyz6WjYe5hY6wRGMR
kBQKP7N30SqAIEApabI5uIIAnScMmSReBzHaHYfC1K+WnZ7J0VUSvZ1F1E+G3KO3surhwAQsZkDT
ZI6B+RKRAEpxkbA88j27lgy3xbSMigtUuVW2+DrZYSyD7m8g429Uckllz/1zRJYGZQhOYQmRd+Ne
4K1Tltuy31x0CsF4L3Toe1bYOdTwOLqJzByN/9je/ODy/SWWwSJX0HyzbR04SiPEv0tiJmJzs5NX
eXPR7i7uWxtzqhfBWaWpRz/wLz2Fp+VuOZGL6ONdWoNoAIq/wuBZYsPZcbMiyGSytREw+gkPGkUs
F+yui/E8eeltGj9FeEt3uKAcgpkI0BN7iyKltb6lGqSB37ByHy1w+vc20TrnS32TpUBvJUdfZJ2t
Pjfhv41SgcqMy5nTbQJOPtQXcdRPn460kpEE7Xv8dISXjPfJrSBNoLev1E3bAsn4WoDVet64qsjR
zhy5YA2GIdRGj+RC4x3Gu2cP4SjGuAgPaNJma57gYHCEJTuGSONBJZEfTyUJkMg9bQrjmX73Lk1Y
UWSfu1YNthnpmcvmH2l7XBBJMZ4OrKdOiOZjXRx9TEHCtNCTQnzK0IP2vhltosDeTN5VgUbyMHVP
192x2cwuYusSg2A5tFKVZIH3eci1EUTm2uLFYZ9iH+jMiEiZUXBmbvw5BXkoDSMrkOg605P0QDX1
LV9pQs046N7J2jR7PnYuIQPHZGPB0z9L9Rvu1OOGDJnvceHk7RBbbBm5LCE4hFwvJt/Hbtdzfgj8
Wd9GFLAHCC+EBap4JysCSdGJWzdNpqF/cgOhcrSADU6sGkvxibGG1UaWIm+84NqB5CjAFvyCdYoY
4ThXSOXoX+wlbBq6RjZIYqvkb+VuPymy2fuXnh1aivPs2j6oMfpqgSP4CV9vmYbDWZCDxHIKjl8o
h7Iz7KZGXJFRYJ31hmBHS+03jvdrhBisgf8TLL97kM1p2rqnMJHXTuSL26LZZtHKZ/2jrVpSlKrH
f+QwUEvU+hoyWYSgk41kx3IW8oyNxOsrncFjPmP/daUJ5sUxYxo1BNtYAs9vLcgtaI0phXxomEi/
WpvDdrx3D76l6mncXuGc0rhm5d7sju1wurliwFc6Lm8bNRE4lPCHR4yubknr2BTge7onuHG50Zij
IWJ8l1KRFmYuF7fgngDbb7WKJhNEY3t9W19PvDxeKL5UPUYkefn/gsXcwlZy0bdVDhFcjQHcybg2
RDln4jCZEUv4DMcFIXdMDatE+nmuC3h/GMhZizOGTWGsIDvjYWsfzVBPlP4dvtzDbSQMXdAaQhC5
jfFY/3SghMcxdCUJAuGSqgeAgNYInSKQNYftGDe+GFRdpmQQsQ1+ZgiDNO2FyKp1Ij5SkNDSjSEa
bk8ZRpIlDIq1kK/NAlj4LXac4w+lOBC4+BbtZ9NfPVG4p+XLsbqYkoqCXgeAOXPRmAofyLXRfsQ+
qdcWZo4jV+YbxMt9CV8nBSftvyRtViBMkkvRhmh3+w9YmlPXPfrYd7ZxaCUO0GxhfZTEE55wIjX4
/GFUibEQTdIt8KHrZQvmBO8wKb0D9PSTY8SrpNiYJLkjEdDebWrICifNSzkCorIRtWq0K7QfDxa6
chcCkh9M57AMTucjQVVsVlB5SP+fUS/cgNtr6qVfkA84ycwggZ2t5y7aOkSjolpmEtB1f+uWYoQ+
QDZxEvfn24229TXw1tTum9a6xG4Wqqez7jTH9vXuHuue5aalvmjsO4H8WQY9LO5Du92F13ZJErEl
S7Lm+a+WcPpetrSQ8s5GnQ5sGvXonJbwGQdYjJ/lgUutyta9A/X6hdrgyaBhLK/Z8FrtLSXpmJ9N
VswxT5/IGrg/+7mgvj+JWftuEvlMYirFCQu69iPF09tIhpCl1iSVvX+Uv1qRDgG9PdKeKKxv41B1
1k+KMlmKdG1X/CpB8qBD9+id9wMBRSyJCwcsGIj5M3SbD1DfxG+p65gDHpOmce6SaDsXpGfQKU4p
bXrBCg/npcyP2K/LhemQkW8Kn9Ywt3FZySW8PVDs6ORnogap/T34ihRT87HSKy2boOF6SFpzjHut
L0n0ZqtCu7uL+UGEamNbqhJtu5iQ8goU0UK7axZVA3/qavQ6gmt6+dfu13HjmBwB/AVx2iVyZxY6
xMzFxiwaylOoFNoSD63wTJ9Y9D8AvN4ySjlLXbxe8zR86SIIZ0HV5Qbtst//FLN4az7sGpEYXZbI
cqLoKGH6YvekphxxjuQgMlYfor0afyLSZQfSt2M1Yn4/m14X40Nl1qVhK17NWsu4K0ZXURiFp1fK
62qnf3NEtRTzT/JeBfSwdpITXUm31MPsBUbOCXjDPWrqfIsCa5KbyYZeOWMdvBjHl/L/yfgDMC0T
0qB7eDH0dVw5AIJJ/JYVpggt1d5ZOkA08PcuvLsKsybo4V06NK3VYgVdFKZ4GREvj+ze33D+UEKl
7AhZVukZJeXhnXpQlTx24YkvRjKrTV6n4VD9+vcs9GqAJFj8pKU3qyu3RR6JcA7NlFBdpBVZBAZ/
BVw2njLGdv6PUtZfp0NjQVe5w9VqodZWmsktCLkwsqK1disfjw0PBlzBHSemE7pY1HwHSae1iXr/
+3Oly4RzT9YpytB2ljC/IbIbXFUB4KRKRnbrAMOOcuEFEA5HJUGD+XDNimR12szLiojkdcF7i30c
fmUAWRPY8EOnHz09QYria1d8R5L2fO3vxEiN6I5lFu5146tMj6LwR4DJJC0u82BJAFNE5UqMGX8i
nX1uRtznC8DR56i+5BQ4O5knYni/CL3T/m66gUhv4IQduX2szwRAPVUsE3qpIUFhoD/xRkc+2Pzk
pDgfR56kqYHstQOBzGX22jQLeI1Q+MvKAGC4WEmJfHgs+a8iA0f/PBPnbUVA3u2GVOZQeJY7eTst
cdVB3SDUH7b9upPTPsr+SzK152I2JQY6OT5a9YFVQ8Z1sGlB+QdhncpTWJ/U4Hlwu34uXEK6UZyu
i5Pmb7L/r4/TDDgi4l7M//bC6p/mDXndpk6/oxMO9zRGSmmzLw4JMuMSfz9Mx7rxLSkY/lHhDteV
SI1FjW40dyauLqoM/FmAzfR0oHx23LTZQlDgKRPlzsApOfgfaSBu9GUYJ8V/hDE76YVIrOQ8p9F2
uFRvNtie8cDePOpyXnFuZNxTLQ9PjkWF2FucHY6ROj+gcmUttvW/qJStzHGmBEft3ZaNIWDq2587
CfXiT4PR+ooJZDkIQtZwXoKaHY2lrCzsJ7eOK/BsOxvmcHSRfw/qRJ7UGr+oHCgZqViT2fyEnlwF
AsmGUprS4S4HBnLzOKxDv3qwVFPD5GbFB9uZKreaGAx3ZVcnX0IUj3UB8gS5d2JBBrOt4uVGhXhY
GxElr/R0ZAYd0xsIIVMxQWfX4aaDZ7nJzZqf9YJM3tkTDTrfTJPmR77b4hWCZ68AxfwwuycHvOmJ
VErEAHxttS1pFdMCcN6phAAaXdzC+fRhNhE9AtDSsWn4bDIdFcMvm6fC/sL9nnaxLZmu27/DDQvQ
1InglyPiheoZh8W277MUgTnVhd0JbjovmrEAIlzxm/aw3e4+DFAxJHsV4f/AvhzdH/wUw3t1int8
ei1aLalUgAi5Mii8GDcPfCdJnvJVXS5ugXVn2nUQeJ1GuJ7MBu6D4Q3iK9IgdStltwtpGzDFC6EK
fUfrwpaKC5hwqM+hSNYKio89eqbsdBkxiNyJFLefOoJ7FjDcPUe27+TdGw9hAaoOyMiAZzaKr1gD
fCrmeCtugfaAPm/96breYhl8Rn235XxePb8/ovKSaf7Gd5M1DKtiWoktQjFK4XNmWQkp+QcFoK1U
Xo/5KRUAccTz2z69qjdWO2B4JOMdf4ksbNeyGFI4iMEqr6orkSgSgCiZCp5zoKIZqykvaMBOGBfp
uMtNf0fzQh7tcmgmtAhfcmIfkmmZpue+jSft2jTRFoJHlivdOr5j+L1g1s3pPiHled5bJvQ3seFa
QDhxJlDL0aHso2Vih3/9dZhUEtzGkmnMxXK/xPUPRLoGtPz0igFDDAc2+sl6fBXCLQLud6eA0gEr
txEX1/WSCxuroO+hzJ4KTHR1n9fuCkfSnXVUGDeHIc/mOMnO/a9TXj8JN7Kj2A/mN1ZM2fanCzxK
NJ0SYM+bysNoMUyQDgAqBXfGzRZuQjfJF9vFJSot9Wu4Jjhp7/B+dFZzuFyTsFDnn2GaFuwUTX+x
cuzTBVeXk7qRu/S8buPWuq5YLtdiSNjCRSwyTeBGfiucXFETAA6FvnD9gQjnIcM5TeixyPYwcbGJ
3BNPTxt5J4PpYVh/OPORIYSlYY7bjih2tmlX/Lzusgq78Px/rChw2lrftao0wPI7Odl6Kx9YgzrC
tOjzxjHyvE0A3pgUdsd4BPe/cryHMlmyPUTqGgpVHOq19bYyx/KW1GSqZMPxvAezJDQ8o29LJAZM
z65yhmDtHNv6KsKmr/HL9CSYn62DZl0zxR10MFlxGhZ9wG6V482pK0uIVVFAptLGuRTV2tGwzIpU
yClqJgEfTkEzPJv5XF2kAPmZ8mpfJXaKcU61uLowAYoIPzXu7fu15r0hIMvhkFmmeuwtS68P+1iK
BQxifw6cuwrTl/VoAS4Lb3zMrRDmpaHd6RCHPGbTvAhv52bWOqEx9xbeYK1YMmfO7aUXSxRWn21S
xvpbtHaS1ddoCz+/AyIcqeSef6qFmNKrGNK3BZCOVPZvduCODRRgnINEySk6mBTMX8DL+fxO8GBg
AgOLGEk5g/2yDzUUQIUNMtaIvzd5PI1il9YB5nTrXDnXJelpHr6EScVQ05AGZMrbkmnnIDmG9IOT
v4Fuip20JzOqpTbqGvzqhcmDd80bhocpNzTvA5pXokFhMyiLCCN+VdYm1x9L766H9owOeMfvG+VB
KGumahHjLtbjdYWzqwaOXqu93oJ9Ry8Us1GybxJ29gvMKxYwoITCb2hA2hHnNiQkKyUdXTa6+c6n
HHRxSFf1Ucro2EH75VqbTy7eBw0nf1nEro4YUnzUj1b7X1/VgOcGwAuIPQCZtUfaWvUJhYJY09R2
8wonxOwiTqfs2DkDU5pUXro0SecVzffJQkRfDLzWydB8HEZrZTInYGnQ+oMShfbctOnJII7NVHyS
pJ/WGS8yz5VuS/JdeVZjlaioByp7R74qxyXQF/NTnbb5Yn+X0kVuI31yMccKK05l3/ZFM4NIPKl3
/8+JjvHoQ8WCFh6ax8edcuXZEQKOSjYNVWfvPVqUmwJ9UkExkDyPFUwfX46wlaKOsG5m1+wm9i7C
P1uHe082SxXhFzdmlt1fC2wIfu/E0vR7qoPYye2gaHs1CZBFaBVI2fx6CCPS3C8ikkquugrqjSFO
YFFU1NhfEACEmyaeymSmg+fBkx6k33TI0OUWvtVeEFoccfhuoUIahQWqEx3gXe3rfQ3wRES2gKaw
rwzFIEgLnA2/GNatvRHt35jZnPewLN9ZsUFLUgn5nv0gpG61Q+wj32h8+cePHLgRfJf8qVHnDXxG
+H74nsCJTT2+AgOWzNFtt4BIk3jSwjufk4g0QOCG+0mpQZI44c/ZfKKvSR2x/mfRdTmSRx4FyHLp
v2GsS8KOO6T6IlSnb8c97fZDWJzeuFZXiw9g4haexuceqKHMLrbKbYRrwP0CE5HZU3H6916SpJC0
Vu4lqrYjfAtlgiRhihrbvcYDVPr29vkICZznWl7H7vIJ8CGQ8tmYuqQvoVLL2sK4BlUZF6nyuWoT
ubuW2766ks38E9g5r1dkOcKYHlI6z8eVTRVfVqp8AIgtfBXRPIh24b3ZEO+jHslKuiT4u65oVAl7
5XrPKvrHWrtmMoNxBnN4vDRMWnVeKVB9Bb+nCXDE2YvO3WRuk5u4sAbU0meQQx1hy1jHUUxFl4m1
KnfsYYjJgi4zY7bU+9/9Fej6Bh5mORL0KwSCFR1JUmvFnCK+IaUwAXngoybv2RQ7BqpzZtNkOXxc
XjEwW2ZWyuaFAsMHYsAIv8BGEpyUIHerPiwFHaG67pwXfZaqBwtCaLbyseW2VXp8X8KuRkS4VHgV
eEaAptJ7liNAF1pFd3mChrSIuTCD9ECRVXQuhctKPDDxkdCW+zB15IRnC+akFChEond28E/dN6c7
Kg4aSC1neg28n1BmISdQmLy+Y0wRrGj23zACCUO9zuLjIuNKNx9UygbErsErUWxxZ326vujG0Psu
TZcRfy9hJnrls6/VfT1LF3DX7jav59jUAN4U637QU5ncyn9nlZAIwVlt0QVR6RjxxAdIeV78lQiR
x9NUscmRatkDVnV75JHRnPes0Kbf1xAeOHDEwiWIovaskcGjifwNl59ePBCKSq7eOlJVxm3AACXy
WyOdP+GE8htUWv+AQwO2snD3e0McHLM9I1k6rN2o4IpZLtwVEuayBOD2tmqbd84ODJhOFnhSYFs8
fMW4pMgau/TprsJrBqPeQoNk7G3wsD0Uk/WSmFXOY7pQkEG8fdGvTHvwURMe3JqnTZrAfSWks6B/
gEPfGkO11ysjQiqC2w2DgqEopG8mSDYwLRluho9u/yP+5fXmgYA7U/ASP5Efa1n9HMtyHufkkmpZ
2piYDo1rfkWrmx+tYQme8Bsjci9Oy4g9duJ0jtrVdLiUECitHi7qYB4sx8yZyvfqeumw77CTjJ7f
Tyz5je/vi4QX9AauaI8cpWuQhUw0XH/QB2zCpBTXyukgGVx9xOKxjslgi+DRcXqezq4z/FF8CCzS
rx1YnGsRKkuMxgXReKLzbrEBC70IBnbDjwH1bGZaaaAQ2W5ACyT8VPCwsH73qI4DLY2WzJx01oJg
g+WWSf/tKeuwwsXzxpt51fpkIUV6lwrVpkPx/OX8QzOaeM9gHUVRuwH8mkw49SHZmPUPJRo1x/2q
vVrGcdZueC/OQT74ubkS2/v79E1kjea3tz4QqSqlpu6fwhd7fYyR4SM0GZypobf8NKNZpoD9PTI7
C6EUnCfKJjli2OOly2IrBvu8og6knltXQJejd0cvtOYD2duc0hozfliNyVZa5wkE0WUtewJpX2jr
i6WQwZaEnc/3SsKTB6BC4fAnw+8183sI9VQDasKoHfk94HH5NGoOcujtLv/SjRNiIYVP52RzH7bI
p8iHqXO9Nl5lZ1DoP3L2tSIIQcU10+vFq9bwHah1RA9MfMdWbYkSrIxPUHKVT60uPAvxeXuOPJ2H
93J8Zdi3lL4d0Oj+fImaca3cLZIIGvVH5j8BgkvJxkFeYPmHSzuwyFQp8vtKUsKyo0z2rWDtTcze
BUL1quHdSZPfKaPsboB/Hgl9nWhjtzjYT8ofCDzNQG4PY7F7+xf7kUr75kwilxsCMe8x4VxsV53i
7ponGyfxKgx4b1W6K+xkOFhxtDq6fEqFUIcNSJiXa+L9pEXYV/7KRpu3PQKA6u6LLLQRKU/kwLbR
3KxDJg5c/t5g0XCptZJXd5C518jaGWjcjkWIgLeHG05pmtWAYHyc4iLdxx83g6WxNYSiT6ONq+ui
f57ZBQZ86KachBiHNlbkeOwls/RGX3MQAc24RjqFSYA/imKORrN+iNEqJNQaAtdE5iDYasz+WvQm
38rR2AuOO29gIuR7BYxcCAylOMxz6AWeZYXMsC5rnWP3CWSEm4N7Qi5mkn4e1GDvwTrhmb5Ay7xT
jYjZRXqevNP9SOi57vrkot1LLHCUu1HHejKLmdVCk/n0A+nDaxMSNEArHBV+JZlNZQVC2vWun2zt
Tmghc/krtV55pjIbbIWNBQnpe5MrwXsWEgK0uZsShz8kpqk4EE4jCwTjJCLuIj8Q33r6J/Ghllz7
9evMFpRg8Kwe9Ni3VSdyX/StzBttTsVruaBQLpDUG7Q/qmE4e+zUO7qfWZbu5OIgf+cMWLGz0rqw
NQ28xkvlzVTNebUuQOxwV1DEul+9WY4vYXH3wzb6KusPHfbm/G2HX1rDas0k8yvcMaxUmqYWm3/u
asSaV8PIz4eln8/YFFKtCz5NpexuODvg03R3CHyPMBLQIjUs5KeIfz82O8PO2BH4BIrR41C2X1gp
IjElIlVLVlIM/TRWYym2lR4LR+xmEqG1G7T7RcTCsZASRLIYAeqXeDVKRE1MHBjoPmCjr59y0zSI
67nBMzibNBvxkWnzm0Ks8AwfovcCP2xsc6LGlu9f8eiziUskz2q+ftGDdKuOh3zf2KEj2gW3NLcK
+hh+lcJkfltZvLdnEEouN820ByTsBL06VD+dv8UQjc3coAWLj0V8EVepNlXK1/+Ps2WR2st+WzAO
sEDo9Co0ACfUfC7yV8jOBidYX1esGqg7c442KcES9WF3/LyY3t9uU8oo+0D31JL/3yhH0V9JYp1H
LH7NK0/lwvWvh8fDrUrdpUmwKH2iMs3dlt9vYNkzXOyakill0mznu4QsTvgdgNNHIX1lc9VdcQGg
NsOMVk7rZKuJ8i3ERvFej6QzXdKbm7mGCNDXrPhfXnf4+BsllU/nGQDPHJv0C3giRotBUqCLnoBr
qKIv3/FDvhEbOTp3LPiPKpMQTdx1XMFPzrziVBN3T14N85P6J0MuSNfaMf7SfVCmqdLtBKvMIqC0
D0uJdFcWkSQlJO02HOkyn925d/QxFhJkWupWNkxL0xD5TMh7ypQvVA9AGc8Fwy4BuGJc02E19mvi
TI6IfyU4wN4VowY8i6dYOhuC6CwXxOWUHC9BBpLc+lVrosPSI3ccXXdcUcY6uF7aK8yC/CDA6uab
Qx2izpRqM769TIkAu15VyAEmpXrdVR6ZeDmkX7xNToxAAZTpDIGjKQ7hqP5rH/c2x41fH20ybEmB
mMofObAk5VWFWVnJKaWxo5pdb82M5gsNNcINVz1kPC3vsk7ZnHt0UXJcjOhqIh8+C4w7uVZY8gmV
S8+1PsMUyBH/izzgkIXR/fsgVOMIe2KUZNaUKyDmV3ORPNMKFF4eW75yh8fudE5LbrBfg6jaxM8j
45GvFMobKR8k8/UP6U1Ktlydky9telMU2rroSsLn/ZpcjjTxo0Xw1JySkEJfzxmlncccyDsyteSk
HmoRaEU1IH2PZBpFllhU8SlcqdYuWM58aLqzKI97lLn4VahPl+3Z+jQLF/CEY1eUTcxKWyhddKl0
dmeyOqZMMltCK++j+aIYnJI1+3s4DWM7ZrnaSq6HAkbieWwMYdcmUY/8VuBWHMnZcZjFekfQShcM
xLsk4NpiOcqoKv2SueW9BlvViI32blvls82apIWdhW2BLCzBFyGSCaZzKXh7FcrdwMdXIfIs405V
P3Gyb+hOEdbew3eGcfCt0Qfgw8KLqAXJevghcI5AWkisTs52wbB3yuxX2tnMFAwudnDdOv29eT3/
ANQMo2oG3D7o9gfkhIt2WLkY+YNDwVIJJPHN/z4oFQtSCYDdET2u28xhmj+OxaacANh2REzNPXBO
croszdP/Vpgy/H8TXpBl46RF70rCPPxzErV/n4gSXRUzMjPeSHvsxVZilr3BouoFzyOUhO6DhJVb
ROqY+vJyVjymeo0ojELAb+xj2Zfz61EyNrBipZ2DqSvf1pe/kjyShI2fCNiCO1WD9CtZq9+79Gb1
EM34K88eBf7qinmC9HeN4AerFcZlUoOe3cnCbvTO/39Ip6Su4Bl6qAroLB4UJSsg+OsWuP02AIBA
nxxsmYQNWQVb817rmJxZUti/ahPzMbxsvLQWyYFPad0qdJo8qmcdRlmZzoyq16G+6Q6HQGdHQgOt
oX3JO/4YGopf41CJadE6sAMMkswybwm0jI4RphBcRDxrkt1f3puYngOwGGBB9or5y52xPJQp425G
PqLwQqn7nZUXgpq/ayTkMcq+kG7gLw0CejbWuQ1bK6rpVQziHTA0EfGsQGy0zGk0brJliqPDGaQM
voFqexnGmtgUv8ryTJVhV4VKJbk8UEI8dV8iiA7HqeQHp6dA0WzO5zmisUIR2IBOLS1rkszQll8K
Nb9jmECBHq/xmBiQU9b2H5A8KboFmwPDF5QrD3UV+H0cIbcTjE1/Wa1LjXCowy4x+NtP9YGJvh+I
4AZypjLJeb7nF2DftBGZ49XBuETy7peyYbk4FUFOIgdTd66wi5I5ms8yFyUPgKjoXya8qKb81+Ct
lixjtKTHOMskF6o9lyYB+s0xqiPSRfKeO/aIX7JI8CQWro0TKyilqEvdjL/HTWEdlbBrBUiUecpm
DDMnXneBP71MZjKDL6gzh4sWeAKfPqr4Pc+4nDSh2fkU/oglm1+D6mZEEkzFtioyAgg4n3aTyBFW
1m7yRuLXvv2XRwXEuccXU24Ez8Vvapy1yVOk/TlnRuMU2x7qITbhIPW168bnkZPH8gBPdsucZ1Wu
8NpM3nDZC7RSxe/EYSFyUEqD8ZBwmChAsBC7+rKxwl7/p/48t+8FPu5QcWMZGuyhadkASxCs64Mq
7S6Dq3gRZ08nzUdgFsC168BUdz9ZsisIkAG+6W+KFD3ihl1MrnKMR9sNKFK7Jmsiz/OAqg/qHwff
gckP8pDomOEpF93QJHYOtuCQbhlCF5a3qU22upv1bGh36XIN+x0/9eZzg7uLoO2JDGAIk+asCOSG
MuU2/8tSuQWdL7Zg7qXmKlemhlm59pP8FCLAe1Sqpou5/g2CH7ojod8UsUxfZBb+DGSsB1Wq3N6L
9zt1voe2t1xu16tyR/1GqEftdeURy2eDNCmfBBUF2NOtEPApT/bZ8vP1eCxIBM9wT2IbBxyUQUZe
BUMPDnFtjqjgVcXMXGz+jg8jLTWtFvUWWPWcW7Dov0nOW4Tg5hCXW3xHTLaGuytZL6MCff32mSZZ
V9PRGbixZsublw1NJyqSXRbKQVWKhpaOcmHc1xTnHwW66UtKCZAlWvPiAmpLVadjOqub6H5lTY1c
CBL/dL+PrGNZHrcL19g0Q/zCndy4sP6LcJ9D2NsJhXnGb6PL/HNJZvezFkxsZgVJIEkmENZKlVT1
OW4LNWUAqigvKggo47hP+xygLYw5ifUgsPodczAtVyKZN/3eNKHTLDN6Pf5NkYjuQqcNU/5YdNtv
I/oSddcrdbz/9R9urTh5fDzmiENvPty/w72M6h+jd6sQmvTMgBa49gqfxNPsfqjPzSqCcKJzgh3u
Ks+sbxwhUkrG/Rlh+4YISs9MKJ2PpKq5m/Guf1NsjFUYHo+fqY4nLgKtVLuPMB8SlX03pTFm5QeT
lhB/SXUk1ZLWZ8UDTRKJ84vqIUNoQGYenc+KDrRxSB+4gA14C6PU+tmxFLU0UULqPSCJb6U8qiZH
UErsQXhwuMkq5/0Ugs/hsbKP8ZDnTb5qGQ01owJek/a0NTK0Nwf8h1jhLidZ+q/rDETek8d2TLIP
VcVczFcMQBG+UXSM6iFrll3W9mColJPjdJhdSnX+uxXUG9sEyikXWDdYEz42XdZgPCg+QmB/cqxm
GmHeAl9n8fm3IPkDc53/0FtfI7mPqA4hP0BXS7H3CoV3uwPC8mYBn8Ixq2dF7ob6DiycO5NdM0w4
RlRkUNCnuoPdGuJXv7+B/bGckgbGRW5W8VzvWAe/OHHoWrHgD4qUk/EhLCQT0jrFG1VHISiVZ1L1
PFLCWNU5cT6SxNjEBSh6+sBU1NiwJHhhArm/ANg0kWt8vdLD4IsczxwqhSY4cF4pR0Pa9hcAYssf
qyjfcQp0fAtC7y52DApvJaNs5H7Hwys2EVduDYuEHoY5VXH7ftgBM09EC9LhhZVJNylSxHmjJlow
ZiQuvQh+/WKk91kDPNZWxsDMfc62R5YMiIhnn7Nk9MdxRRP9+h4uZW8I2Zy3dssPEo6xHL6fNJbV
emfKfY695szDFfEWTJ5uZCgCWDCAx4d64eCJHcOUpcpcKUIp3rayzU7uZVGX3Y9xkw0o5nqmXuQQ
e0m1TTn2HTQJQRo1a+Uf42cf5pavWGhOUZsXjqX7z373kxX0Vl1DtbsRPcHAhQKS7uRmNALJ4nmr
4Qa9cWNALNFspO7WOHdmG1AlmTES+erIO1Zgk8saWyptfZ8q27KbKkepZYTC9CNwhGqREft/VhzX
psquKsx14uKUATP1j8MnwbItmbnNJNP5n6cqFO/DiNmBkDx6srk8C7omEob6FY5Sbs7sLO5A7zJb
EUsg+C0ub6CwqgWQSnsudrbG4Df6jhbQAQ01VMA5AdrW2IdEzgz9aV3Moq21JvctgfywrDUXV1Y7
idHc+JTbGBimfmP/4gAl8GRhwZRunZwMWvcwUXHRiKO5NsXWPxJFokPNJ3upD5np6EWLD1yKN8Bu
E0BSyLqiClYNrLywQytysZxe7kqLdi+9ESvPEM43+EaMTYiyyzYSTaowtCQDoWtVNVZDYOf0nO2o
7Jj+VsZTXedGa4jH5kwW7kFHIlSKAo4w992YmbmTpzbg1covNW9k0tJhloBKcDrBQKS+GZGPO5BK
Nsqt8ej54rSO80Tn9rLafbdMavfF9CwiNTuht/BA6saXCEzc0lnBulnC7XnpxiCe6JhMy4jJkrZ2
A6a0xkv0S2nlxOV96FWXMLv3jOv2RkEClYvirh08A2vt+EESR+FYikJ3SVL2RB2/L47LZBxUnSci
OUpmTJOAY8mMFbQykmo0aWNCrIOdsO29egQ5DDYrZpgAGuCzIZhq5b/Q79/nLCMeTjmXJMfD6MmL
R3RugD4WCgWzGx28I+7ksRXYwMNzNBKUV4Z6yzu2gTXX1LurzzhmPhubym8Ix89cIESKhgLGnZ7o
ztbH40Nb0IyDNlMoOfvHXwWZ2QyF9ng7BCGwdz3vfcAu/y8/b6pH8nVD6JbyEfn2fdmLR+Igfw5k
RfAnSlMbSJ+EZ+qwsYskXmDtnHuIgFc3jI9c3M82bEvUX/zWdvBFbSUzEE4JiWakifCmRQhiipD1
LUOCcSeRr2YnLW7jvjm4lEbET+MUFR1vhI5jLszYq+u4LrFtXwf6wi5cQeryCllmDufC4Q/M+4t+
LrdL+X6tzaKWisAMjDodkaHkF9P7JMuAOklRLJzL3GLxPnqjSpF7t4hDLt9YA8dFX+8JyxRAoeuK
nvifI3sxTdRSq7MqaE66iweg2AXxYTd/cZvbCBMevRwRRdisB1Ta6bvJ/o+MCgDGJKE8Tk3RF81f
Vo+jHLBMPn4mglejaVllNxdkExMHXZ9xmEhLlI62D4R0wQMEVbTskkHLOjKKUyyrsOFYhdJAbo4V
QhSruNHYiSH9Fc8vj/WT672NcBES8iTAw/HJZ2TnKMOxZzysN2FWpQOEOH13gmtxp/ZUZk7otRia
nV5jCAprT+niz4p4BW5jGio+uamhYnt5fnMeS1i5CUXVF7f1li8o8Pq0QWocq7HaLGgrNDmjjV6I
38MIEU58k/Nlw0qhL/5Jj//OUOcGdIeArOb2ZIKCEWe97+wkFip3QZfj/R9LUFH2rnFhh+h5a3GG
oeej66VzbN3nhUd84KRJU1ObnMZYHG/YU5TM3kgClFci7ZGQKpHOxqKS/YmWvB4ypvASUco8ftGW
ZwejwvGsvss58vezGKh+sq8IIZDsej+n9FFyTXCb0A+qYJdL6Cvj5PEAURdlfR7pkub00axz4Rmj
9MpMp+Y1+ZWkM4rw/pmMS3V3AjFNfM9fBzSlOzAhjL5q6a+wADIln+zhZucjKlWuyr3jTNVLJjMb
ZFlVzrrSzDWqw7hQ7IgoNMM2z+5Ns6Inm6pwNQ6psYxMVlXDc+qBnvzT7hYEfYwd5wecUR+UWi9A
gK0mEqXXApfwqHllUoLYsC7cI0qz023Z6NZOhSt7U2oALw4buUV/vF4Q6JIMtBOLkB1HV1slDRqd
6+qvz0fJC30tJywnWWgvCOGn6Agzi1H9v3S6c/81WNE4Yfw/tISlr/FD7iNWIfZzGAFO8GlE1ajy
DuRk1SNRaS+i38Et1rHRy4TpDbhHIl8P2Z4zxYumb4+eKxn/pQrKY7XmSTAPhbzB9d0ke9gkjV8P
jT1bkPpX/6eSrPrzUEU9gBPomHg+aP4/mSDFCMHa7C35If8ra+hZgNB2x3ExgI1kQzEzVjEVmXyg
24yM3XoUXSkPsHdmGMdUtokG3jz8I4H6XUjBvDKzR34Z0nHLkZYU/CvwoIKwNS2yU5O0sk9KFSJ7
dV5eH0RAIc/4eHdPujdXHmSE5Fa6xOSA0axxYiGo31oMs4q7F8utL3WH2dmtlHQqLg6bZBXG9oQH
GDAZU9N+zSLuWgPQqzePCPiCgJKyC4qofSlbA5q+FkVSAD2hg4i5JFJKLV24dSMnLOdnHeWaJoqA
4hwmeJqKbly/eRhQIBifi1WuOrKQS3KxI7iQD1GjJsNJJXz+Ytk3D5fw24ftsygDXekHyhWG/Cwm
efGWF4RCjUd60cschB6LwMKMFH6N2PHw230lKnSW4zik8ML3VVCC0AAFR8qzhrAmMEYwXd+fkIhI
jbihJAu1/GloTL+0goAr4i5sf/+MfMosRRjrsVQdPosfZdpioVfx+IUh0lSSKtCw4Ak82WpjFdI/
QpdDlfRvricsOG7T3xMYZA5x1Eo2dz0yPaBOlhvGcCL0XHoSNRQBiRirvbrKNImsWC+MhyQnhYe2
SFP7FXJRvFRvicd10rnhDVeAyOvtLK0EJbL3m1nxfF4OkBVWac1+A6XzteMCe+N5vmv1nLWhoBUJ
BnE8z2uRK2QQhF6NfzafOtsRSgk+wrM6hz+o0eylYelUxZI48ASsF+ayTpAcwJ7lnudfLRhGT3ee
H54umRm2Dn7ZSDMulODTIdNkPnxlcsIKDS3lq/Ul/3DWN90Wf5kfbvd/K3TVMKa+pB3gJdHOx7kN
b93raGhqUPbWL3T+scin9ltbES/ocSzd+iAnrilneDgjg3tQfIoULcAsMFLniDL0dSVji6V7WFiG
Kcig+2BlRLuibhEs5TJU7cbM7SWtF668GUev8mkqm76ynQAu2q4WMWjaEBiFX8RRMUbHrIV1zKz2
shEM1PojcZP9rYaDqOdkOtA73Ucdd/3ty8HSaQs1GW0JJR5OIZ3cJwosOY+rLaMAHQB4hWutBwSH
ZTpxTcLXtSW97pQXQTmHXIHIR52ZQb85EPVekkSKfa/BfgD2rpXeGYR6acZR/NeGgNMlWd81PnXp
yjiGSiME5NvuuQ6CYtWeWzkc8JKyp04c97bOByETkqBNXCHZ0lxRQmycxWp/urMfAZ5Ylqp6ONtp
Q9NkXnhJo6HVVvd4XZthHB5lmKZT+CPUdfvDc4tC2Lck8o6pHPKX2voZp5NB/HwuYGIRC5spxhtD
+068PoLI0Zgx4NkPW2AFCJPgLewOHcCwCImLbi3U8kzUdcndQP5HNDtf3VJ2QWmhkAgBkzZ5a03m
YUJiu4KzDNuOXf/QWjK8D1J6qa+tDxUix/f6FhD21OYCpdudUXkkZ8pzgpQ1tZCJVF9XrRlw+mGA
lTZz9eu6B/NfUtxieX5mbawcUKKFWya9Fhc7pwj6oO7pJOizCWNrg+7fNHVwnu+iH3z9oKh2oU6O
2OUcpHKlt22gjRl1y1VM9g711Hc1CTb8YPadeCbrEBZsutArdOq3LOud9XmiEN1IeNii7hLMgC1Z
dFgxKO+qh6Asfvv8j2tJP/c/zY91Bi01ikSOGUMmhJM6f8yHlRpFpYARJjyHkIeltu4TqYFQ/q69
O3usPXbVuPd6DVULlEk5h4zsqp9NmcA/JmzSvRjrXafZcKw4KPZb4uSp6xMlyv0J/krKs4vc3ASv
YCzl7ZTHIkWphdyvQb3EVwrxVBoi5RR1jmu2+lyQHOZPHTrsQJb3cc1X7i9ZtVXT7kj+vtzq1AJp
Nj//pS7by41xsaiJcqjSih12pKJR6wUXw6agFZTjTWV/8WQGBHyZqKocjh9f9Kq1ijTfobNlfWo9
vDX8y/aip3ieLPkK/j0PA0lFP7s3R1laz4CVBsDnkohaZ6w0StScbtOABxf25wuBgvAl77Knsd2F
Lh6thPlid7Xc+M3/JswYczKiyHuDvpU8DSAeaOO4B23MtFj6H1jE+YXkO3ZD/w/7mYWTpgqrCvAU
qVIhs5GNQWRVI10K2adpSq2rE0zfIGAz1HWdLJGhs4uRGer5yvEUoZQGz11ECRYHO+8yYhAKEtBz
kU2s8B8xUUcGB8jKwrqSc4xiVYSY2VHap5o9WpFUQFGdiLdhG+nOewWDQZ3VVeXdaC08Jbp7weyC
QDtTRl4iYgVQEaf6NoQ5NaD0rHk+EvVap4zj8piB1zojAqRllzB5WdC2hXPIoCg6EOb8VB2oD2/j
rT7mME5oPjT4gcUH9hwYrk+FfTKnI0ncFMtKBuXcCeQg9sZOxdzMW/23oM5imwwTmYZdZuK1HPKR
ncT/kCUXMnvZDXnJ2A6Oph9fW+logEkYZke+l/7Kc3FAq6DsxRvdqxkFuuF9j13mrPZSpsiXxIrG
KHRc9Y7skLaJGxeqddD4whtCn9I0Qhm6h0lCFbcoCgjgi2CaMDkp2HCrL8YYM/VnW0f0NAgF9Ikd
7c9xWFdiZpATwUHLwQs7jQJvDrgDRLwdkS1/34vFiuksLu8PeZrLGBIs27ykiz2Q959lwZ5KVzmf
ql/p4jDg1f/NdQ5hsy6B3Nn1NyfqV4rNMgOuKoj7r3SP0esVHtQTe2k2yV/Yw5TRODEgO859082q
JmPPXisY+FF1hK4NvgOXQ2bIheYjhnQTenLOiqId8uOALHMuUYKFzmGPJrUTgJXR8bB/o5+rZVh9
73ATLcy3PhiECFWmRxo3y6Ux9LEmChGR2A1uVKUYJhj3MRGbk4EdQ/bkn+FVo51Zw+lu1IznFxNQ
xerNQNaNMrhNyvcFB7LFQkGaF4fC9jETIAeM2Va/pIS2C+XpQ7p5eDjcekuz7osqXA6ov5U+dZ1B
bi5b5cxNm7yaEgXrgcQl/rONaugVo+JI4kbblbFea+BF1LRZk1cg2NHHzxa75Gz6fadmtZ0jrnY6
67IYJmKsdxQElxX8j5w3cXZaukef22mqQO1ImjHK1aTUUJcHUY46//TiDP6DyL2ZA+jH2uy24p0K
8ny/dmmXEBjZ1ZJ/w+5xYgIrzPZtP4HY4VzjpxuVUBNeHKtsenLqJrbFZ+AhkfaUEPfdr/8OFcKi
W0h+Hg7dm27uMdJ826MgTI23jJVMhnoVhpCpuUaHbChSHHEfGpbO7Xpnj2xQHDZ0ZOX2ul7PJ5yn
yNVBgNbEeEET3/766xpW7ddTw12Es8B+ww5pgBf+mn/zcTcVbdbflLOk88qmCrUjImbxT6exJQ/p
yI71X38WfglFfKCKUgi5wATS/oQnbqR7VUDJIepvfTlesbCixkfFuatl9KIzbXBV4mVXvOjkhFTm
NIBBht3nsgUZuKslM88ZdOARAh5J2pjcCCLyo/0x17fBWiJskCtxiIinfh+qNIc4Wp4TCfjuKWQp
JEq05FZjT0HNIfMaTt/o2zilMyp5msQ1pxbwAr4z+ARnkaM7vvffGXA53SQ68PeJpbir0pLT+8xS
xTM3Jh2q6hEm5kvQcwT8toczshTtLxGXm1RSwLApvfaXzfigEXtElHofZD9g8wcS0Ht+wMAYMfqw
oi9O54f1o8q1sBBy/m+7IDzyCd+KQdD4dQsymlnhvXJNhXehj4IUFKQ8WVsxOiViuQ5oYWd2wzpR
I+KNqDc617nOH+bMVVbb8aMJ1cWpUdamMUAXC2xsBh75hLlZkMPL9CpvUNmPgusDusT5IwLyBew1
aSX7MITIRbWoXNVZSkD2e0AB6LEiqxYFESg6CW9/IEVBxJ+yH707bY1P2g3AjsjrEMRg8H9toWi8
K4DRAKWRXaqZX9+ymU5FupLVneZqLlglPdSdmTKI/P54cOEPd6ogSm24FCa+34Qk/WyGOco2XHvR
cR/Yb07DprIJc+bh+eGjGUj7XTykasdbQrLOttJF4r2/BYIfuUTwFsAOxDH6m0egIcAvrvkejA4L
QVVHhc58pvB0sjXqXVC0etHBqgHhWzfmZfM8sr+qB530CZP1xunV2eMZ08HdL9q++nSfYSerY5LH
XwQGV0MXAahRKdvluZoax8rEZyy9zFG0uDFhVPzTIMstasNfafCQPyxVzn5QOWrR2BYhhwkhRzvH
wio1y34Y+bWe5wj34u9NX0/8+PK5/X0//3onmudTjVTFyswUvJ6SG0ZdFS3E7T6JNYFDQL8G80hK
0RypSOkxLXozFdxps590ghugLbnEl3myxCbVlJCkn0i5Qdxxqq+8D4/gKYY1kbCjM0+X5DkreUbN
p31HOLoCkkOWqgk58WyjHeYAqykO00TOeCLUOZADsQzfovRDDzddjt6Zf+haskOf/X6XLnQfC5da
JkLnNMnzhihftSxggNuNIKngq10wbcv34HHSyxolOdSUbmiGnjYETjmMEBT82AJQwOUj/VdVO2/j
ynM2ekJhhKO/RiycL+ejSjDAawiARzrAtOW4dIgFZyKOUICju7u8KdH+rMnQR9ehTUogg4sZ5PCX
EWwkdTit1WpApK76yRaRETErR8BKYgsQRtd6TPQp2kRfWmtcvIyaKRMfV8BQpqA3HKoQ8kiPZ8hA
7942OreIVV8NDhxRvYiWWDi9CIesbHDn2kT0s9WyqygjShWOLq3LjkUZH+IiiAbUwXRBSsYJKEaR
grkjjpGNF9PKrGDPtPtk14KkazF4vC3qVbnzL+zbr/n3uk/NWGajFtDV1lcjLJw4lVAob7cFEYJ4
C+s/mYz94f1FqY99PZoNP592eBw83Ed5UucYQnhE67BIPGYYShridQvCSqQiEUSK++9+qTt0HZto
sdDWKma/vZ5Ed2uc3jK5Jugqs3ZAbxeabEXRBeQsnSHYKRi7p0+7cJFgW1fyZ10PS2LQdi644iIn
zRczgFLDIQytQ5iOxUElTeOGPrddXoo5213Hgha1MmgY2caGwTQ3bZWoAPo6XtSf//JqGrCCEqHn
hQwWm1tX246nkAaPPpkTLHF/ljPnjdgZwsAvYg9LzqD7FbAj7tECccg5qwao9yAGFTlqJ2AbensR
GhElXTqqOUJ/C6hyac1qdXp1laqwZQ7VP09mRyBX/1iVhPyY3QmnTY9cAsuMerixm3sQGceN6W+J
JeoKQtY/2+kcx9+Wz2b7hkShv1jyy0LukLK0jTIMKKaVSazEVQDeysVPvFXHVEEavXY0ApEJZWun
OvgYno4I2fJ8lBeWOQpcmI2GcRJzOlDYRI27bl/KF/lRudG3fTwjoqALROaoR2tXiqHPd8uMxQVW
Mvvr8mmGtBazuOC8e64Qm7JEToxYgnbHQ63WE78L7vnz/hnbbIRc9dzDbYE3xzbn9vNtFDUaDZ56
kBoEXVuZpgTjERAAZ7bv5/l8YR+gdh7eYVoeNg36M+5i4KvQOWeDMqLmYtiKPlur19K+ovQrcoC/
QnLwiDfnm9oHLYJ19B+Uwxa3E9DX11xpG//YeYoCw3FEBY7ieUu/W3B3l3ozle0ePvDfyXdOKWkb
TED2+LmG+OyI2bSfD4cJWSDu58AvYsZdYxeqeTh2s5scAuZlA5sEq8Bu9kfuK+FyLwvE0vJF7VFL
m0kHSHyaJKpp1JFECS+usyqEwZqTPSnuxqEFYvhemM5EByy2cwGZuD3Z1JgeU9wp6cRuPnIheqDR
OmhN4ZuyOpeMbWeDrRs7wMgTkJgfmXbZAe3sGYKuLrDZC5XzfrRxdafuG2mNBu11D/n8MyONCrmp
Rd+Spdmr8lL1kFL/le2hzQ99TExLl4rNUbVLYPkdPeWe6yOKmnRV7wey2Kz9HM8cupBKgTmzOAoK
LJ2xIudH5Wk5Xa6mj5vlvpsnYVr8lmEvIyrbb+juznZUpYMgfWzerdD5SGEdYh1xqPFxmgoDj19V
SpSJDYYRhNRelY1RggxEi8GYD1LUuWlrDDTFf2p7vZlSmpVJnfIuROebtTeBT6ILtY2c0u4qaGGc
frXxYAzvuPvEFu+/k8cSnoGOg9XcajRh+umF/bePiFhHkTYfbSBmfjO+ahKPbtWFvqGmCPv6As+G
Wi7EBeX7VX/Sbev1mt3gzGTyQl7gNZpCMs7OMud+sBomsrrEWVnccexNI8R6GMTJ8XHQ61Ybnqw3
IkgKRLfB6UwiTtTPOPrqrerjMgYFu0td23o5a0KBRDRnKf54nKd3AOGfjVbsGcS9V7YhLcnPpOt3
Kc66ybxO0euyOJuXXeGCbUce2GG9KPOs8DSl1g3dwhUfEYHQA4T0WVA536Apu4ZE+KWzaAnV2fM7
VQAiD3DgRwZ1b7T9Pqp66Z6kkXi23g3eCAhQ0DdF6ZnNjRxL7snbriZozqENnxnhFf1917lJwlYb
vtPldEaljJe/+DUvJDnN9zU/J9ZTH1rdEMrxYjL2lcz0H4k14mbTr9/keQNoygFech9nO8CA6W+t
FYUG8lHmnibDmywqnldTnX/wrrMUK2DB+spy7PXc2hNGApkj+4BoeWLhT/Tn76LLUwhfoLUO39CZ
tQUmq+QTxswad5JBpK+ACoy3WWnnzhWeFUMVkFy4K2JnGgKirDRcYqVo5R8zYAnbjjX5K6aEuUcg
X9iah2sYWhjDGylsB6EfWnZCx9QUjyFab/9vHUx4Ov6N9MYCiO0WfcLzcd5mMk70fHA99tqklaUW
K1ijyKEJlh79JcTh9gQgIFEMK6csGFZ9Ul0No4ehgOmn/2t+GwqLKp7di3HzkHS+yyK+QKa5QceE
uX2f3aV9K4JAqJqOs979j18i8vm5XQE0Hs54KvcAwqwvU+qDVbMxxfJfqcD+ZbeHuTy3J8KKsxRz
MjoiLQtOQ0Ype8UyVFR/fX04iNgHb9ArkDoTuzijuSalwoNjFxyGsHA7HE/zi56QXm/HUVB3Npi7
r3Ny3zoiONO4dSfR9t11R0IkuUM6OGO+relTwTyUcUSbkRdFMw0Vn8gs2lJQWlQUE0vy5Ff9W6vB
fyId02vQ4dZLI8bPcZx9v0pwNicZrizQ1eUjT94DorSH4BJ+PTGcEZ1w4aKh455qFeOdnHB/sLlD
IkL/4hPQvfETcvDTueVCp2L9L1A684K4Jp/FahvSwDjusMBU4/VT2W/GPgfM77it5E0v1mB4feaT
88SumLaSKmC6EJn92XrVUvIyZ0gJoEQnddacjze+QUzCF5nDkpAJtUwop5gA2J9I+1+MP3YP6ICZ
LEf/8ra+zVlnvK8kQgzIFCq6antvgOtobRS/V26ZUrWVqXBMwf2SShwJnZbnU3KzKnl8IzEQRzry
u6MH9+XIdSLQN8gBKG2ZivFGbvyORX/ulShyrGs8XilkSLtr35HoSwQZFzE5skKSZaDAggNUbzuV
VnXNe8Q6gr3Xbo5825hMCKRqTP7M5vzeNG59xeRxvnQbLRO9COfrZ+saDYYgsypAKJywGvgYmAd0
iN9vL/p14TBoxBgG2Qm+DszvqSlDmXJZHluTatB4My62/hYXhkZyXDks0fwxln9mf/pZ1hmCcK9w
YRadNvVNDsRefotl5rJqG425G9MJcojTw9+K0ftKnf0P+fRK16gVzt5BLYXqxRb1EKTpXKxY0fDo
fKJftjzILCOnjAZkFVbh+yYt+jMh+F2e6zWbWP4SGbBK5Pw4Bou9+5SowY7Z+nVo5fB59MmflVoc
G0kRG+5I2JDIwKFqSVHlnIP0D+DLIHLbvEfF/arFNXpua4TXl80MSVHBA3/GG+9++lhy3luwGpMM
SFTffolh0uh6zdOoAQGYJJPiXadH3bC5DCp5FkYJYieJYhgO5Q0JGcF9dsvVLRW2xvOrYY2sgS2R
B0JKBTc0aQarMxFpgZgLcq4PBsCHBP1iwmdOg0vLPNlp9vrOyJCSAODP0VaRfD0X/ju4kmoK7D6Y
c+IjCPS2xjh2M7xIh8/AUewrNX8IO02l12DBu5pweOoNhjRf9fWiiX6jyZGkeCmy6vSmnabufuIM
WvO1LP0NsNrYHcpBPDMJBgFS1PHLamK7M6f7sO7uBaszwapGbF/pH94WPNa15pzkQedt+gsOPz6y
HCkIY/wEVNP0EEgb0zN/R2DhZ4AucGyQNHL1ErmqcEbJHz22RZQMDT5iC224bnVz9dFpOM8YfIUj
T+a7R9CKENdjYiWpuDn+lptdBlFmN1pcyZ61HRVce2e8Ud5TbmWpehH0pY8JlZ41+ZeJL6M/WhQ3
mR4ngtDKVHdx4aBpErdcMCp3r/0lD1uXG8KwWoeyUawpkKn8+zoRsGdBKf9W722Vu2rv7eh7hX69
47qYtXIxRf5k8qG2k2MVxIB6GcROmVOvnQ86Jypb/jMj0dtkYSW9jrYpady+d+YPIAMjYLctCi7C
vqPul4SV3iOtrZ8ROb4WGzGPd0ehV60e4W94q29UUZ1OAfLeGtrxhwVpbuRFnltVDaixNJlofyDt
P/Zbw9ofgJl6doolO1A2o1F+X1L6hwyfGPDV0KkSs/kVVX9QLp+nwZ6jE4LqQXOyDEVEBp/5sAL/
cqlWPXHnemRYn0Eopoy8g1Pw5EmOGvp6oEQbEAxa2GIkCUv08UbPqs5uU8N/yZnQNrk4FBWByYXk
pJOhymUoqXkzvOvSaJDiqzGwH7TQm3DVIW1ihQuLoFehqB9537LXW6CSimjM9DPDUl2riUu9Ss0X
ui2TTz37jl05JtOpmOm9bKML2JOjNKmwou5vfQ03k2CDRS7HYH0sTNmxgYksidTYSj8DUtryvE/a
I5WePzTPAkZs/zGh9LYst5nrbhEwETqND7Z7+OsEvp57K4dRwmJHCfn9yk+owT2CkpJXSwM8MRnV
TS381OZu3UOMUdlk+k8sBOibXd/dVZ8SXTp5EGz406vQFPF7nSK0WV/876nnoFuFA7p+6U4H+T8N
PeATzWNAeVwAaS4y7vnwiAmWz44iMFrq7by63Q4YMqsF/duYVI97k3+R/6Sfm6o5oDczxdg4whhQ
Lt1jQGuldmKfjnnVLOW6kCzkuFD0D4x2XjtiU89d9xKeaPj0JCwjPHsnBmBnYf18QTgwQaV0QAxb
jusYoYfmjxuwOA0NQliLPCqPdBqXsA+8uAOKX+ddwhWwe+4IqbRdeAyIynmzKMexjcvFJS4SHE9m
V9FFy+gdI0/kLLthYTH8bqoNLfAh4FMce71Llpz2pchTTVmhCRa1qDeHTX52riUXv61KRHTdzfll
i7fz0LVcygms/DYtUJ9ik+Jb6hv0tOBzb98NWDF58bdfYB1R2l5GIOjSGH/ZpXFkLgasLxs63cT9
UCmxV0msY1AKoVw3uNAne+NeKL0g1q6vCFmEhEhDJXMzQwZLBlx/rcEkI9SvGNNWcyZg0bGHZUtl
PsCLV69dP48mKeSwcF28Vnha8syAdPSHELDlwpNg2bqs8493UeY3CAroGK1Uu+i0gyn5fqCMwrTk
AiItZ0TqCng7rAyTxw/EaZagtLFRihaOZgDQrB3UIF3avAvz2ReUdGQLoaW1E0RJUuFNhVsTypT6
ml54eCVoYfUxpufb3gvTS9xrK7sxGinfBhrfO9FiPxKxcOsZBV9V21E3Ab2DvjhNv80UWWUSXJVz
9poVshYqtWI9luyI2aSL/7yrSAzz+i/5tX6uGkv3keUa8l16ivyx9/YBPlWjQ506CUD7OQs5OQ1x
VMQQfbHPYCGgZd5FDCkzbO3qaOxsj5yW5Tk0ZBpF2VelBTZA06s89+q7TZwVs5DSWVvRy+sTOU36
naJg20JUxnLRbCUiMepLO25wtFLZYUDxfeBe7vHxVNKtQ4rF23/st47R5Les/lz3ClcUBqUvASEx
y52fp0ey+fpfcxpy9gMksDlK71DHJ77VF/5AVjBysuU4MMZXf5U/R7zj8RnvNSAKXLtjhv+KUD2U
+FOZUOdTt38AKAFb0RPpIDrD+3JdeenLuQ+Jz+EkVRvQEgTSCfBDlBElfQ4iyY8oZvTiymeMNzYv
X1rFd6px/hSSuy2khkEQfEtb9uJIl9uHw9LAcjnmbyUJTju7d1UfywqsS7fodaLVl03yFsXr31pw
kNcnqOLmAsXv5vGopGFBsKAcu2z0+3ByDYZlJKdpLn52+mjhvlizl8IUiTtNxjwNFzjvLAjaBmHr
9sP2geIdPV8yO/Bpx2/5A/8Ar1bJyrXKzNbVKBlpbcMlXnZJHtC8KCzik66i6dIL/OubsotTRxte
Mc7TDhc+TuvRXI8REIdVec9/Y8RhYHDwdrHnjcDLE6VgVSajBtIbPVvgy03EoVEH+mYTooL/Mg93
FBEudzdXUmTtHjoI6YA/Zqyfx02OsKEsvxpitnikJGSHQqCXBrlPjKiFCKAguSOFU5xX2O0Ei7se
QM1vIMhkknSn2e3nDHXI/R3/MDwN29RoMd399Oh1M24lmMKAnfiI64HWAJHL0slYVswEPi1QM/1q
4G6RP0mYOOMoNSmCbSs0bgsOZa2VR2+JwMRc0Shb8CdZtzk4CbCSxmBoBnPCflqupjzAg8llqqhX
K9/gfKxJXR6tdLEfjkH0TG24wDrNnpTWPiM/o06sxXAm6djV5LV/BIx57jTi6gMjxatv9n8hDZ3a
nmHZbM6B3lqz9n50msgF7otKe0KcGrq9JCkTxEC+dE3tOgR0JyHZMnSJOQq+ra39QHlevP10Jl3D
YFo8r9Ky0rhUHRMv8wY9RYfUVDFy1ACJHK/Fd/kD0uTDivISxOum0OkBqmmJSru/9WiICTK3JL0e
p4usvV3fh3HR0wmA9OIxPuvHn1fXIO1rzGQS48OnwsCS7x2pXJwJ1ue0qNYXkfYj6U9e1sNff7O/
PPhNfo4djzLua0FZg1rvUHyz9lJPJjlJVmIG4ROt4ZyDjA8dMdz9+9eWOW6xqhlKbkqbWo08Bq4b
qgnQbc0w44b4SBc9I7IK6Q9S/fNfjxExxtYXiN469vytb2Zb+H+WFgEw25SmCbrzVS28sUELOW4L
q4bapAX4JkdZ8GfVJRpruRHucL+As2C8mmPo/bL78NUU07oCxVrA7gRCAn+F9E7pMTeFAecIRPxl
FcTACCgkxeiVd0C4hX88hYBxL1f5K4GxrzAv8XRUzeW9Iwu8cjagpptr02e3AclL4eBBtSvP+IB4
Tc/xC96dFE0wA3tu5mcB5F+/oyO8vEXPCnn+jIlranVjgZXl5Fszhz2gGQswh1XOqmA/Tu8w079D
WKNtZYs0eP++y5f+yB9t3hsKuGp3kt1Ol3kThAmtP+QlLM8zEcMFHCOyKGcaMog8/JYY+6lzGZXl
nYfDX6JJUEbHWtPJWv8RWXNLaB+76TA1fWANWh3vWh3v+s7BPUvLsqEB3g2EYI0wRX1/HSY5dGyg
H61tPdNn2N7hWIPgDK6jItV77ZCVisBT9nOMdIM56pIbUNbWNRcprbXIY25Ad7cUpZ3F9cjWzFJe
KDwJwE9PykseyonCApTZhdqj5Ofnjfomxmj9b0Oo3N8SeBJ/5y2njTH6Ge6yuMqbg40SJGMxaMmE
1eJyRlRoGzqjNEsB6bow6Y9hF4Fep6I8Ct9n9iNVJzSfLPomQiBIAJE60E41iggy3LvvxlZQwMTa
Vy3I9r5Z1m2Qg22VZusCXMBXbn6AQZOEWoAxP/0lNomPvnfDKRH300BQzmQKMMZnmPxOQbgec+Iv
VQlLXZzTpya4viSSFVNvpASHbvlo58xhG6cuVcsD0oIz9RUI8r1h/Z9Zm6hXrKTigJtPm6FVZ56D
yd1VQJtl7JNS28AknyhDCol/Pr2SHmj8WGmbEOxyiCm/nkDIyLqqvUf37Z5uGTV50z8I6otFnkNt
13QwWYNC6t3SaaQ5NBO4Hd0JRUJb5Rh7Lq1AFE0cVryGEIg7yaYzUOot1B79RHIELpaLJtXy9lx3
KVAMsYKCLGfT4ycWnV7eDVCnWQ6JfNkse3jRROySNgaqjk3zixOUnxxI22T0Ky1DoiFMuHHmLV4F
klbfXsFiJADr3BHIczvQChanOjjMXAvGxy176ACurCKARiyvgvTKLy5XqRtp8ZiCPFbw2Iytx7iW
FqY6AOXCYdOQq0sArSTw9fe+6ur9NE2OZ42Z/qn1z8VFj1a16ntvyB3y9Ntx+s9aow2VB4EfhORV
oFuJdpOfUlXBKaF1R9fnpAW1NVHLYzVgmv7xCqmsb+5XOymKvUWFCIWmcjXfIL0d8dVr1B5X4Mvw
mApZbJPIYNkr4MKq5BhSZeLEiK+6jEzZzaWNXcikDFa5iX8YVvIgACsaRcJrkcQF7bEy4r6n8Wq/
qwiv3ZIWiaAjPG3dT4mUSUJTthNIz3aFWcpmYeB9tMYAxa7PDMelMWE0EYhGXuNRgn0B1TeLZHjo
SCf/LnMkmoa2/set0fI87+ecvqhgrpmeHyzm3RteaBJPrPXG6ty/dHvbQdBqlcETu4Qi5x2uI/qw
fpp093bMXqxJa6FfSe3plqYuu8XoIf59YkUwcgw7yOeMTG02HcoIua88oRWTE2fpqIYjVemOvCEV
8EEA/b9RjHuBmrcuttAIl2cJR6HwwXRljTcYFHqtfUz95lqBlTETuhESN/nvrncEcQwROdhPlJ/6
rZAnl1a1gHx9gypNpNVcvCgGS2xwwcSSQ9l0ZI1CTZKYxj+1+YQ8uUByoDf+I0AfmEszfAzo/q4C
zOCp1vGRznTb9oRrnELxkybc3Bq/9tTYsV8FxAP/7IoYOTvQ1mdaHy5nAquDIlgWHhDk3o+rqipV
f5Gmf8zpWWYONYeict3UZafRsQMK1whX9NK9mO2SfMqBlV9EO2m1Fb2NEfW4wNkFSJ1NQUR9K8WW
ZelFOACIlLhI/joxBxZBjrQM/1I5olLY69I7PxRkGFlZHnJuoRs+g4LpPuhyjQrcUDuA95hmrf30
u/1+bY6cYGxVq9HrqBmgZyQc3vS+Zrr4zgKVas9uUKjsCWdwJaRzCb2GsqpNTLA2JykxdKxG2JnI
HAfvJULowuO7qcGw3z98rlTylkcojKuf61Wox7nxk6OT20xsbtlOxgtXdc2c8d+IZCTOpBAl3WBk
nsa5da8HcDJftQUQnZEfln2gM/B9Psa0Fnk93LdUs6uVtkXm4UUDcVQYwfUm41pCdcrBFFr6IqJD
UODCZAJKFcSRSlvB8oZm2avO5IELAIQ67qqe3++/GSIez2nurWJQXmq0O1SbEAtQmU6Y2sSOxaGh
sYnpowBMkWnxAEvibzTFMLZanRjFZsRKXrx00b/PC2GNGb835vlhyOsm/l3DKWLLtEhBLAyZHN4L
98Y5bKoCSMqSHv8BTKX3mdCfzSYij4YO5K9WDqOb+aCLBgaKGwrTNPKXY+LJkT/ruMI2yfVwo1wQ
qMQ5WcjKshNhictnMiZM5dNTvM6BfYndOg6Et06WZZb3v1HYxi4TbAxuM2+TSXJ2hZYm2MU43Toj
5Ti+mH0z4nQ/Vcb6dFbgTThq1ac3cOuDDG2C5NUmlRJf6gvT67tVxWf8SlolEOR/CdM6QMDF6uRW
QLheDzZoeS1+m9RHfqmAMzXd/pO/2Dnd78aYRuWaYKN9RTKh8y5YNE3qTASJD49mcK2xGUUB4385
GkvvsS2LSZUyTBcISOXCdB5GVg2FqQZ6EbnTveCofY6PT2uzmdiT1RnrRTy2CkhxfbWPoBIYfsEC
4dBEhid5MEFuNYCHx6kY9fFrmDzf3fXKnEWhQotXXF2KHiZDiM5wSJjJmYhr3052sKNhpi2vxtPX
V7uKJQpxWnk98oqUcsYKmVf8Xp53yhkUVg6YSGm93NCVUjZ0YPuEyrpOJZ/ks3m6v974Dsu5JwA/
QO1lTGWqgoOS2fUsFS9A0zOo67ZC6aXZpmp/FXJg3MM9hgFHmlnG2gnsiE8c0iGdd7xvn0iIlgOc
42cYc1t+vpFIQsPRkRat573+Mi/Dr6JggIpo9sJw3Rc/dDloXn+vY8j4ymsRoQdQfv2tpWwGJWQc
K5JG0R5Tpr+diyktBbqU1FC1iks9mzxMHs3CX6iZL/vt+UVlo16a2sO1XeFHaVZoNP9yV+waYkCf
qH46C+QwBA+PUXewj2JelFOg+ApI8BIn0dmXCfm7atLzVJyaQr7EbpGTtjrqcGGd1rbqYQ2MjcIZ
w/Orq85SaeC6LHWQSgcRvw9rcooddTz0EEOhbzjjXxDJFV9lotqFvU+pXqmsL37rrdphKztsMIBE
2JKY78EORGzTSxN0dgrXFYCc9MXXYj2B54IGHzsL18+qQu+0Mxbn8oGBy3PtHZbt5K7yoA3psKGy
5RWaupsqMCFsnTHSN9JRJXAotmil4CC7jKja7l7tqhhIqHw5VMO1e3HIxub09ZSm6m1obKLNiZJr
d0o5F6tvI/rWEuReXRZ1N48FFV78Sc5lF8VLUOw5rqWtqY87xFp95rwi8mJnKmK7ZwFbtxiYS892
UFovAVHQkmrElLdddcXCSui4DHhEGA8sbLjiKFKgt2aNIXmcxNA8ebRwVtzOjjMFq5HvQxaTTylA
kbjuOpBMEMCBiNJF20C6KhTmEOM2R6Yd1VwpIdrapLeBd8h7vGd+ZaoiNRjmS4QQOkV579q17j59
IMkN+xwE4nvfTcD3aYdfvajoysNcIjRREGJiT/W4loGoUZlkx3JoPZo4sLjJAEjX9g9zY0dC+G4s
J6VK4ylTx5zJIM6AjSVYwj6/yJE6/KVA/FbVHqDHPrn0d1Bv5GVTIwnsbPRr9jWcE9BBZ6IhN6R1
c300EeiM+NgzOjjSkQ2u+lOFINaMDrMOck3TPTc4qfMDF6o3Khv5s85TJjuu3ShyvE5i3CwUA0UJ
ouRvL6HLClMjv9hFS8iNp4WPnL7ja981wd1/WAik9HZ7SywuuA6xs5GPpO3Bdj+WfhlDK74VXlUs
5gnuQKXiw07VtbNj+zdCTVKPqDo74YpzGwwXrfDUaV9454ElHEBTRFXY28Cqgf4X5DccniXT/NU3
WNcmp/F5s1oa5BZp1+1vwQhSeA6mcbYCe1AIpFUcc9YyItwEmJ/G3CGmQ5qPJhoaJpF4BqnkWp+W
dikS33wfIkWnSDn/Z0PCrCeErgGXWEvBXKYGFKxx8/ViASlg/pNtS68wQ6yLWARTu4rT90JJWukN
sz9enfF5i6v3f5mY5mfLtCu59rtxSWhvZPZfktBVXKSPI5x0UUDDEKc+2Xw/y9suytjWoKWnAtw6
D3l40rHK6QMOMCC9jxma20AJMBYDPsuGHOUO88xJMJk5//0+QC3/pN+5H36oJYYo+0h6OzNatKNE
BPalftjLlCZGDy8pp/tALNEFmUsqGgAdnU0T2JxrMiqCHq8oKNh7ZhOvcp9ijijZtoz5skcQAe6y
7MrXd9r1kEwsATsZNEM71BbywQHoImoXsf6bqFY/vSz7fkwIOITFqTsVyzxEcuW/6HwMkCCkMIYi
kConDaV9GyymAz/NkcKpL5789EjhW+lhME1Jy4iXiffRyF/AeaeocF/vCaUbQ6vkv+0QQkFFDckg
FTvcAj84Dpei+UwPzv+9LIhBGUTwawhfX6jP24BVKBfH01f1ZprmZv4oVtFRW6asTegzm9P9YNlZ
TSv82efKpL+nL148ZZxn688pHDAsbq3+TJ/ks2TmmH6EKGkNYHBmywT+/tP7b41ig9sE72bh2L68
tycJ2Dh+CyEWL6sWm451PD9yg/U0i4bbOx9rEbGMiOWO3THm7MdvhqE/gj9u+jn9xzBD/kJvJ//P
1Vi+WFLRmflAwTnSAk5jBku+yc4U4yPpidGuKLjH84vEgGQmgloSlu+eForwUaWg8cTxJRYtOqzI
g+7t5YDFiiVFP3n5+UlIXYT2fGG5cHfD0g74t+m9zD1uYUT5qjxShqzKd3+tBt5p1p1UOlXPCyFB
5QhOWPw5s/V8lHOjpsHgfi8iwi3/Jq64YOpRqDC8HU9PwDc3vHWrOnb12cSge4KMIpiYiDaOs4j9
Ic1pWG2mf0nOZTbWiXaGUx2ViwCI38x5ox29rzdPwO5vbe9NfALtQsMDmtntgkDuDyUvkluoepbN
tlRXaoO6PnCKo8U3VGokqnNPmgMQnMVlb6FHRYGTaXfgMOHxeC7SEgtFjWpPhm668OmOdfKlCEZF
obr+tF4cuRvMIKZyMQxi8hZzjLZevQhp8rHsL25O3KYs95CEqqAhgXAcRdTDoOF1BVMj2ys5Q34K
DUzp99BPWXtmoKzcEkY7juO+/957zg7+MnmormzClWnYG1Mx8Zj/+VN3E5ZE/4ewD5/mOcRPwsYX
hSNAJY8bXl6BCkBNPcEkwU3PSMw5B+t9Qrsf8SZP+cKbt6ZvNDcaA6q6PHjuULe4TkffB1Jf7X3J
Z8GyH9FChz8snNQT7DDCsZMru+vFukUfDNY/7VI/qfEP3VKExX1gdQ5GAdT+s7FOlrh/Q4GmAf+q
uovMjuwmNcPSWc9lg//g1OYVf/7zV/4M5XN+27nBU5KkpppdFZ/7eHZFZsMtktB4fkR18QSzIa/V
n8DdoI1wPGDtffqdRIitUOM1FU/jq6dk0FGAYvcYSmCghZFJ5ndegeOv6gc8nyXksQsepFf1Kgo2
fQurNCDacnWyJ0e2kN+Lpv5IlaBslrx2VWuDd3KhpGZuZyqA89s+57vciVxMpn7kmdlibUaS9ZD+
jyCDttXXvpzbVKzyQPjFdOr9PpS+VPrPg1VbKzn8slMvew918KhooNzcYC5za2reLII0n6IIhZTw
7vFurgTouEEo6OYWFk+8CIWQpmuOJpCDepAnrK0SyFa6BGva+PQgwNJGTA3MlD32aHEgMzAWLMtV
gViQ/mh1FEvBjixpNitvkkVfIPZ1Itu/A9CGtA67aLJgqNNlZifDIpBiS07rmEC8GUP4zYRHvM2M
w35Re1nxdB6x7eqleN+UhUD2skDeHJ2EwT4J72Q5tstvV1fIUn2bhzKvHbHh3iG80SAs9xNhRJlX
X+hb0pX7Y5b4UQPpbDp/ozrSarWOpCLF2YJekr+SQTmGuiPISGXXW5uc8k1cqQpLRXuHE1AnD+rY
sCkqR5sIyIopMpkmrhV5bxXRgtqECrxq8Fcaxz6tarGZbpYJCOFbtVgsstRgjWvpjfNBNGmRst70
Et90HdTHK9FoClbnAOJnjcHeIHbWC0vE6t8h77UAJ+gjtXlM2FisgM8ORiKHwr1F/CRX0KUor/wV
lxOK+IQM48xBU05DURATglcz41V6maw0EdJnyfP2fuUaR4NdWbKpxR5g/8wozZx4xoufrxK8Ku9n
53iRHir0GnSXChvRHSX2hiV1aS53HCgxny9+1UBllKDacvN9rcLOgYzIxogug6A4vFCwt7YNQqro
uby0cAlupSydWneMQ4Tw/H/JmuMyA3knYfGZRVNI5cWTwpWJ0vJLRyG0jSOisdYu5P9j9Wr6Wx3X
2+VDH/RHXoLvTvjsW56Gq+diydaleSjXEv43G5JBL8K68a7llwDEyRagxH0T/cTJ5zn+9LyPOXOm
nq2NKcPvbkWZHRVZz8jTPHQgwtifQkWK/XoOqHkOkc7DCUllYit1g2DdtrDq59NqIm3prniUVM4a
4YWcEwPiD18yDCPocguIbx4+U9Eu92gJJMx65laLMiBUAZOXfIFd2JR6TYpOkCHx/8Pu7M2TFo/7
mqkPKhtbUnfVraZmsm26N1kWKfD3+DpVMJJPvZ6eNVLOpWkiD7KHbFN2yTc7M0yUq/AiTfEHjdBF
IJGsl24L7wZYaYF5mPiXxkR5HXvwDv0S4bcXqCxyGZmoKAkycwPLIrxCXfuFrFy4C0YknKoryPu1
P+l77I/4jf+bRFeT10Kx072WzuE5bwCR/IPfTDNgX5FX9SyogHUNIafxwltv+BFHQzLoRxvrkdVH
Xj/cnHPaX5tppHHFUWA4G2gn5hVzeH8WrvBcnPW4tKFYAhsAsfd5/L0PgYcKBYaYCtoCOcO0jvy7
dGMxVLlSAPBP+3MJZMeuAy2LKz4U3JH4lGOTL3sExVaF7aUu0UZMffpPGZYtYSe9tFBPAg03SWvV
hvMNiZVcrDGlV3Z47+PjZwxP+BzQSYZmQansENjdPfRZUEKdigPcXhz+8mR6Zs/iJCA58wEF/zNf
K1+5BXqcbDhIiSqySxfzm/H6znFpQWWhUfp84v69KLDXxkuSh9cFrsFFX5D2c2Y7/BmnPm0rDsNW
BZeDo82+TsLO5d1YPu9Dwpa3x/uH2B1jDjUWg41Y6xd9M6TAEDFjqufVs2EkIgN2oep/QGLn/Uz5
3DM6UwQWGdQdtpTaOwSns62j4JCUQgxd6BWTRStoflxKxEhQhYv1g1Z8KXiSVPkF4+44TYeEy/ZC
Y+o5JPjwG/BU3um4W9nU9vQwRa1IZwidEnz9LivnEHLiA5DBG6Q+EDMmDalBSUmv9Yo8U4Y8Emkh
4s3pA4u4XGdgLKrz7VYzrKO5+bvcVdxRSQ6k6wg4O8dXFkGIi9XZ7AG+7voz6e/qfpFnr0T56QO6
76HsT8Dpy7SmHMKoBEafStIqGtFZKiFygb7D4s9UKG7faiRWWtyKfm+cO+mxEYvPLWgZ01C83bbB
rQ4ugy4+92RGy04fxizlGvsW4TQ1/Zlz5mwu88N6XX75194om8YmiZVJczddKQeAGX4WM77Fiv33
cEztCoWnUMHd/QOVSSRLxJpuIiaeek4V+0ZL1YxrNqYejm4KUitlHlfKuccPXNti8XxrwKXCHn4Y
J44X9LXix+DvFSnN/0f+rGEKm/xX+IxuHmj8HKfJ4NEyf6+Gr2jtdUKVtWW50jqAKg42HkPmPar4
zmj4574bYxCpmys1pIeHzSQjrOq4V4+wf76MvFLkhBpxBYoGlSudw1TKiDMmEtzYJ3F/Y5MAm7PS
c0JK7SPRXlTMrRFDIulv7uGCmPnikvFUQgAYRomhmGzCwJjVdn3OqQ1w6gIBw+vgrWxO0InCWF7x
BcXfn9PRqlQQxAETFTzUuU4eJYIvUgLeHxfeC2izHVlvYwLnAmQwtF1mM1ZpJTke3NZjNLMwWlww
eEm5yTVszepRzXMe/6f2gsApuH6PXPxmTCsHRAmRscJmgTDVP7/cT6p9qWVaaAHmmYaba9uGLdiR
gRnguT3/NpN6lfO4Gj33pWVMV28YJQsM70+nh6q7/GSA6pj6AcK6IOfen7sCu2SnxvyHN4IOv/Vu
fpVzuU4XLwYOv7jUnZPtqmtUXefpoXAa0md63eeCEpQp4hbuhh3bbmyKlKCqxVyU0vfy5HRqO4KH
f0N1yooh8jf1IdWcdaRqD+sGGVIo7Cz7UzvzwQSSy/DoAjIgnLf2NITT4GGjn8fv3EfkRH5Sy+qW
ZyMBTJS+Mme4NzTSCGKwGqVnOVDH/nYIo7KjMhbmGdVN46gqSRCRcRRPfm62BwcAwXdDkZkCHn69
BSDF2hmc9KFIw5ZXPxSFLqcNPoknSA0IHfgvsR1e/wVFpadaebDMBLvLRAk1RX1UwdSWiAlH/HJ0
nrSwCIRyeep4QX/HwqKk+1rX5d4kqoIE0AhfmiFFmLgzCQIx2ikheVlTpEU80OWYhBW/WF+e8DYH
NNaFFXC0fa7ynuHm9kMv4QV4aJ9vamCypX9lEaKjYJxIvGGi6shAszVRbtnyD6/fEnlbOQGsXZpp
/uyFsej064II5kh7o6SM1R1S7Q+LTiMrWDy9G8bSIk5tsh8WYd5GKLu4jQVu3n8kq7TFKTc7IZaA
iwYPtquQaZtllXwj1cWSfOogImuYQOS1dDXn0A/g9TkocDdXbztNu5AoNx6r5lfKGjnvAXQOezqK
Wwu2gpg/TOqZtLzxqvvvXP4xqr3a4jijYSNUBYPpVEU2ujf0SC8CmiItoaZDcdlW403LI1Q6r5sW
PhvzLXIQadzRyzpQf5kFUY6sPfo/nlahO/CAwSB6j/CcrO8EFjTTsmHXdeqVCobqDQoSfcIlp2rb
ZFrXeHEZnXphbx9p1mIeSx5IdoXzNOXDjerto08nKgumSrdtDVKR7zsYyYkwEBWnBnMrX4GdwXfa
NLEi6M+3cHtg/EDk8KGU2fDSNtcLKk41BZvme2y3lq3Zfo1xXx2qnScivfe9egjkdweRGas3CqOV
qnxFlPAAJsIgF8GYlVLDuJbZxl31tcoR5esNYXwf+he2uvGLNSWB52Cp7bWV8kUeRLcv226CUzeK
k+3wwqroC077QpyH7yD5RS8DTNTndDpKVDqs+36zsjZsoEfQLboTCYETUx9DJiopwpFhzHNg+Hxx
XV5efOfk2M/clPq0eYM/KWmLz2bliijwkuaTRZOail6qyX0I3UQUrPwC2GpuYkILNf5HIc+o2VvU
odWRAZQviW/VStuFTh/B3rRyfkQz43+r57k4hDwfOOKLN7XgyvMOowe6y0OE0CBWfGwmN1TJY0mD
KJPYJbmpnTDJ1KM45vVCGVfEoIIlqg6MOocI6sX3LWgr6FI9hkaqBkRwx806eroXiCVO6kJRXi0d
XGSBoHc/1k3VE3HNBvqG7jHAY2pV60u/v/BFwKXM9JKbSG/TpPfQmw99EBV1yvQqLaB5i6U/dhC6
UEUwJ8qFzNNNHNCzI2912MY0XgC/NAMkcNnBK+p7YxoBta73bdMyGdoBvocYn0aopQ5y+va2GyIh
h+9XYpr02lMW7JlmtAAQFFX4VVWp5TXtVLUtqofnsFRa7ITWR6yKxfC1uVgs4dyH99+gi9h/5HWg
JUWfDuapCBn9/Z9NO0nuD+GnzyqHkxwJoG2QSt0RAh1ShWHCiRKcFeWv/bPSFKQWbu284CgYmApm
o9Zkk/Kha5vcpnf3MIW51Ay8wrHqLUDjrPjLGB3gx5juXelGow6m+2xDOa31RvE1spqRK2TGRNLf
sZLkQKKbW+dlcKLGiJJ/oDV78szgImH5Mn+6pVtZr1iiNU6I8R93Ga1szcaKcb6qi9KCM8GZzxSn
Z+Vu0Ze2hDv2VkSfb0C0a7lnJ8kXkzwTKPYLB0E1IwqdRJLXU3OcsRlEl+r6BkQAXpLHtT3A1siU
bAtER4uV1t2pPjFsy7Si0CpLiIKd1dbYD2ZZs2LKDCNwHJ+u6+giZq6tJJVC555v2HTMhr2cnZkB
OdSb4gHkMmMg42YDW+oBxElzQOt1wfvYMB3yqBdL7BT724zNoy3wFMPR2jU/EJ+VbOVqliFu9tSG
x0LNvuucCzi/T6rbM0N3LKwvI8ZXV9tkm+T6JAXY4h0Se4CiPwXsJovkGUBuJxXd7oKB9oLMBKKI
+YN7UJrtLNZ7vpADPyPWiNGl67wrQdlMpWK35caqlewpZRqGGleEK25pVnhLjGPlOWiyiTbuRQRl
tM1FlFdiXxsLBk+795faQLqvGeDs+UcvVlvJ/s1XRUXE6uDPykQEBsu5f9G2zQC7dhWJm9BQYeuj
Vwskq5lTRgz4fWH6VSuU2YuMHVqOIK423g2S+rkd49cVMmt5ndM+iimNJj73J89hffKapZoYEcHo
kgPnSyWyd1oWvsNNQPHzLBM3OoJc5GQZ9CNEjSGhLFyEwG6yD4zlq6JiTS0xiEIlIgjsni1EMhAL
HVvXfMPdUQOsPdF++alytHn10F0Valjvl/tQMwEWwFmswsUplXqgnd9k09bDp/XlUPTK3cch1KFv
0jizeprt+gUJRMBkMCrpzGdjo5aX23Te0ozNNUo9SoLl/387r0OoHrC+OgorLhNqjzCFDlEvt6G4
/AEJbZrqeYHq6DhGpP9G30LfteseJA8wmTPLSEiYqm34Uj7rA4QhIN3F3T5k1xqcohOxQc/7Zf+N
84uOLE5kW8Q29WDgY2JkIrhLzbB0ri/PI7H0FEZBgm4yp9UhN2VXhrdxPbmkrRKpq7n97/tyDumQ
NLkIhRe94lE2+HHguW7eA2bVq1HrKqE63Lby8eSGPulswu7gi5LulYCg0569kS3w4eO1FqyWAO76
91JfEV+cDiGEVMc1WNDLoDF9q0wodEjJWLIE7lEIWeEC3Xy4205sU9pQ/10PXJqB6fdi4Mmr7IkF
DeQQAscFq+4vCflslxDtLHareR2NNE0cUDrCDKlWXQmcL8BkSQuO8wQyisOTcTZSzP/2Q12czuMg
gWwsqGhT5uybuYm/vDA/ux6YUNYfj7yTbXvKwQtHWWGw1HL8YGlPG6sfg249xl2UGHu5ybUy5RQD
MSoGBlK8JugXkgzP4isL+TXp1zW9j4WGMC9uYBK+5npEJSYoWCQBoj27Y68mRH5b6PWFc/XNzLDt
29rWlqfqnfQLPCBN/TdQ5qeuZ2PprmoKFX7woc39R2n1Z5qgqVd89z/ElSGGZ4X4MeRoW29yA8Nx
HpcwnD6SO/4kQSvh/Mk+YJhKK6G5QDu2tbRHwZJ40PWsLzKwU/QxyGfXKboZtje+cTX9GuOskG8o
mKUbKMKTTkz0wPyVycUzS14E9a8p7VCxTkOFUdVn4Wx9HwQkRYJi3KPGrZ6LVkHS8kO5sdAbtpGz
9tDNCwF8vybTMQL3WAQ5qTHbtEkhcS5V/Kz3ayKuRe1N600xlg9MRset+jzztqEMTfmCisdbLMjW
GrLmVmqygAb1HS+iBfZWl6fHTc7V/sPosMb+OU/cDmVc6Bjp/fETAKVmeq9IQ4JDvLdW+St+wf76
6GfQNzGRX4MR3z9fusGlEJnNwWZBCLSi9pVy1gkgOCP/SUb5yN41Dwy0d5c3agP7PBj1Oh1tSIc6
YYfJ3eyl3FWcYNpwJMeoTWD9EOgt1/JmxTniIbgmSXi3y65Q3qiOvCsZuiHH/FqsZm7xQRQ5hD8d
/KYkvju/BEDHhBF/TitWKFP6RhWQceC1tNzUJEAsOQ0+FDuJS/Gvj2xDjNult0fZMNPG02v7tu+H
ZudYBUViC7WknUMBHLecGntP3NyhuvwCR5lpHXmllvBStqUQIMOCSt6bUxFQ7q+moqMLi7yo3X6D
FwLIYuL0l8PiauPCf5kRKzyuuQHq+NX9qzIKlAiD/0hFTVplhtNYOaAoJt1zA0MRnIYV2E92lg+w
q9TXrfArgofo29QGddZRsQc3fBNd85usGEBFpFOfEAqIs+98RHZSP6oHIsg5Je8WiiRBI+beMA5g
PBSF2pE3CgModzIUKcs6wtOeNVbUzA+qALPwqIb3N8NHF8Ul9tgQdcUR9YB+iXNif2f8r4heVN74
hIGqdQWXXU7iQfaPXrrk/w5rXqSolS31eJiTFY3LKYO2m2ncT08BPyYUB+HYw0KPgLY1lZ5Cp8I7
5FuAXt5B8YBeK7Mc5H54BskBVOsgnT5PjRPL2WD19OsfCDKyRbq6gD/4Ff9FOSy6guHM/pk52Rcw
ZyPuEvPPQEAfQjmE+HrVESI8TSbqmWdeJrXLlHqoFdCjea7pX2EaqLY3IdQxbNFLIvrYU5gkaLPa
vgByQH2bW1O1eLFxBjzHQnEr1nwHgXw0Cu4li7EhVSnGcNrcU+6dERtCfQDsLI0Oo3hTa9+RPtNB
DgxVMfX9qGKXeoyThMOJ1jl3gdtR9S14An0y8Nxyex+dDPArxkrxzpjqt8QVV7+ZDhGzuLYSVSQK
9xfk1o8ceg34xth/2SRYJXCscVkVeZVHH8VPl3T6xgq8elvgVYVfwfFtZSI4Y7lqbGaikUDLzkGJ
6NIqVMaLA2ZIczA/ePC9NKYUZj2NFK9E8NuZYHUSEHDiR4KUQGhmg30aPwsWjZU0455KBbYzgBDf
MJOQhuRmrS5MzBTHQGeugfXN+C9urQGjGpUTegIPxB/klXFd4YRBj4Dd0envBN87eEUmnxV7/1fC
cAYm/q2SnS3Vwdc5eUvQrcnwB1oB3mfL/5D+uYL5oxvlccpVNa++JYBryaCLh7ovFMcrxSuohahZ
x7gNt/+d8DGB2WLvmBiErb7C0YcYtFiw5L7/2E3yiNYBKrrwk6W+qmJPr2gJpiwz0ZCt3jJhlq4c
RMYCZ4vM5x8Hih6mvSy0tBXtidmkqjOQEwP82a2QWX5kcYwMOKOZvRTB6ZLZ5rh3hZJy8jfSsMCn
jFSva9zJ7ZEXE8eUmT6vWSHyLmFcsrwhSfqctzzLCpfvoWHOHgwD82c7Tg/mf+6ZfXbxSl3woWWi
PNv4SlJ0HZYmRhAdcQbforoGq3FCoYEcSl15PuSeRYowTO8etgf54k6401H0W4eHZYO8kEvedLoR
hZHzphasUNqGXuuOJLPGG93jJM+shn1MwaYYzXVGDmOyhlTR5uNIS3o5L8axZQO0pcNI/rzI0xqa
aaQA4YutcaImuKWlQtmv2tJTfcPWoLtxsiB6EU6X6jkqy5sRYJJMJ7Jbyns70luS0qOJSPWaOWwM
gZrYkca1GzGVzLZ788JgWJzIap3se/DPpktZEZgo497boOviR8nvgO6M3AeXt9Pwp0e/wxMWjxQ5
uLelM6RQKWDN/F03KLuBgDlE6wALRiCA5TnMfywi/lRo5woBOQFMLLgFgfhzo+aJfaaTq9AT8xr6
0x5CrDUdn8kphCwLJbfTVFMn2qCSpMTims5hMbeqLtFihG247G5pLHP+TFA/6tAtLeTiRTCyXdAn
jrFNVhZWA5dfOPSRG3yfwr4VEgsnVYXxouHFJ/lBYy3ofqDnAuPLiMEr9TuCUH2amDvaHbc/R1H6
8zo2doUJUHP0xB8Z6iOq4X+amRrs1glWcl5TqUmhU/Oc97gAyizB06FV23zraNS2CiNU5DKXaM/t
tVN5ForyNgf2CjHv+Yx6fH57GTaJnt9VjR8zMlffcDAztzs61LZi1/0w3jVLGQ7BOHhbXWlNZecm
XqGSNStE0svNu0Bxzg8eZiKDlGimM/LluJ3E6fBcVR0prhsLeEwRYzeLSsvIeqNBlD52M2PzOhyN
A9HgsKNW9wCP5bsw5xdCOh9/IGlq6cs5Y+qBS/3cz9dRN9wDMTcjVZhU35J7Nve5rz8+xDczuUQ0
6p6c0eIKRPhmpcqlf7qOYnRbRDoCLInANR3nEQBQqwFE2fKOMlUXHK6e8SigumVQc4ty15XAJ7U8
hzjXMu3LpkPPiw/kL6tcndXHRfI2ry1oykg54oL+ye+mNQT7fXR8saUna3k9icPHcRerTHYaX+7e
e6RL+wVDlxhj3zOdm8iyY+0l2A7leXFqYII7/SZMDRun3ApE3kdFlcbHtvpJ1MQvC0OdZ6nhzMyY
aZc06XBXQ0tP2661dLouFyZvUweqLhqbLn4DXO/8JAbenAroQ5643QaevKP/qW0YetF4TTNu0vpR
IYhat/6GCLkDjp+zjeqGM51Z2Zxp8ftDh1ewOIeXdvvWf0lx499iVjCBuQwx7+wOPENpP6qu7XrD
XnKI4zpJ8Py/9BxjA8CtZxfjQcEEark7U9kpQkvq0v8UFxeCMvPJtL1lbgkPakFIcQK0RfkZisjt
ri8tcQ9wEN5+47IEOGqfBPfaMUJIAyQlDoik+HQzcRxy3j+yx7EJ+qiYf1WwXYImB1J3nzhZHqlF
HSo5LE3eW6GGNoX/TAwVdw3hpLYZO22tAhf1VE2xKhLomMQDXPkkir4lh+B+AIocOvsF51+GOoRa
w8GHzIJWpJ7XIhhtxJgT6qTSO5uhdL0rgptUK0DitL2qb3aIQPPJTZak/TnL/ohIvuZjW01sYkTd
0zSBWdndTVJldWXsSzaqbPzFznivX7Wxexk5veIRQrr83GGWKFmAantCa8skK9pcPE3LVbY78876
KuHRz7xbKnGRD1E0EaXEFOKhqNsgPVhwlUibeSKm1jQnq1ezZ2WisGhsPS4QkHrlpmAjGth+tbo9
kBs6QVbFwMu//eeIcoMxRdk0xsxQknC3m6Uew/wOQb1aTIDGtjyANCld99xhXe5lvkmZghFYtUS5
lG1zofBaT3pP8+g3I9htv7gr6V+XSSAOxgXktDJQBMGvsNUN998rEQWBawG26prIaAAC+fA7uPsA
zSuq+jqm+WhdjUE3h4OaQKDjYesbcVCoHmJn1NNLp96Gha1QjK1qocAthkawGYMHU7tVjqk63huU
Ro34sJlBKTZ95SKMrebmi4jRA4vXg8d2xOreuGjgi7DTTHWutqb8VbyNUHyQEK2R+1+4MsG97i9E
rGw8dZDEgCbQyxFUFNzAiEUzkY54McaZtCOgzyFZh2OWQY4aTkQF7V8rrNWwKlj7bF2mIBPYOGyx
9V/TfrHW3Eo2fto8j9PnPhFPu7VLGFZCGTQS0v/z1F1FNmjl9vklgECXcyieQpTkX73XXuTb+dAq
tvqkQMFTtXkVJC0rr5ykqT/BvAdQbjqY5FxwHjyErm119RD+yJA/jICvHpiDszhzUgx0A2Cm3T0x
fMs3iI/CX2UCXv/ftdhg4oSVZVPRFOnzGnnji3P3FmcBBVh6j8l5kESeFtYp269Q4HMvLzHt2HOa
K++Xcph6fudNnJNL5xSlXNbHAeFagYvyd+1pZjVfV8AcPQtgnpAlnQuaD2hpb2J1QhdJ6U5fpw7D
7kyhQHi22RmbPFMrIenD0t7k6rNui8xR1aa5LoKQDbV0xizFw5X9unDCz3z5ehWIh2jR2PpoHUh5
MUVL5mLpAMfZdv3LnvHa6XP4SyuM7n8Goe+tEErqJRmdzMBi/q85NF9tsuhLKn3FVs2xuOLCqwZ7
NN7CoS+oYYkT9Q7SzmFopUz2kbDFUlimS25U2qyLqQUvyJllD6KGSEFBNSrHdW8AsEwMxlMHNc+q
P/XoB4qPFO/rYMw5jGlK8Fixwx520GzrKOF8btXirTX8YnDRykHKp6+L1cp4pTYcTY3ccj5+xp68
JwVXLZHx9yFGgtdpwTSX9VNHK4T3w1d0K02JErYQ3nEhjiBiRwiNmZio+ZfCUPN1I4l6jC2DbP1Z
AVpfZXSCIi/GipdiSSYN5p3Mk9XB6hOosEGzMKB0gJfR3glQY7I5c0AxFjX4GUnz4iqZgNsZgckI
xuvuIkVFaeIuVjZ4bgCOS0uCsPjROs4Gg0jOkExBlKRG5CT+3R5UGESZdwpQpAm0Hhn4dRXyFsTH
N+JrlEb/UyOyWMw8RnkwdgHMub5bELBbQGMt/9rgnxGXf76VFL8N+EEE4ij5K66yPEvTq6zEiH0s
o1AE96xfci8LXVsQUsC9iDeKbfMoEHcX5QT4jS1mYwL9gkUGixAzTlI2i+kPbm1EA9k0MPCskjJz
p09uUl46JfzCZKqqBSbFmRauAb3/6fYJeTOkXBnexopROXs2uiUN8nNfBqDKDSzya2VDiwFMaghw
XCGb5b+oQJ841mLFTMy8wyQPYsZMMIzFnF4b7iO2obHMWxo+tnAlypW6FpZCsrC6hMHwasRVW/zZ
dwGqWhse6uhZnbru5rtxr9ZLZf8wRHfcoP+/Y1KRcz7pOeYD9RGEu+O4NGNdCtGnRYWzzHLCjxu7
3UBK7J0jyq2nzgZabTPlPkVr3A4GwCXCrdjJAiveKHP/IUhbduDYKLD7WzESEYukKgLvyMxeZI3Z
YAwFg20MwvUl1iavhGrE/Bd+lzTJbfhqooCHsHJ9FW9t64lyo9TelZeyxL3xXTlRBk2Ne8DudzZY
wrUeIf8d10yd++2zoXJnyo9PPSF1scJhYRlYJRi15CP25BurNOjPIlWIxiaSz1RRWMixUmdFFRkA
Lcfayi7WVcxjhM5VFVfhxiqTO/UkKR5fppsyJf6i1RjC5zLdc4kq5KW9m+T7VdnQRCOJKEZ/b9mg
u5Xc1q+iaaHiNEdWriCucKyjqPlLWvzzQY1pxHh7/vP+mV+VKfq8qzKEWFoGXov2V7wsr2wIhvyX
GsUM5Ataku7+6hPjwnYsBbR4ZkrX5AOnRyUZl+kxUNEJMYR3aAhczmi6ZZZe1/HmaZFS1JM6aShS
CEdSZKpM/XGj5kyzpfXmF8JME5mDkDkp2zqnWiM9Yq+AqNu8+7I6woQegFmNMo/mZVdH3H8klYhT
uJeHTcp6Ftu0T4T0DwNPQ0GJw/xIVgYlXNDXq1HaWPe13czDFk79t8fCNGjByBhXnCD6QG8MVHMJ
wNbdc8D0us6nr9jbSnDIhFJ8ucYhp9XjZq3vHVPbf8m0ZvUXBXC9pcoaBWA4KKDfPy1MoyVO9QQV
l4BfoaGLZ/R+MNXfz9b1UCuWSQ8TqQApYUnJvgX21oEdwHwX4Il8yoCGwpSwVetgl0QVE4HIEbqN
VgqSSX/2DGEJkmsDKNY0+hX+6+lKNf04HLygEBW3eLAJklqaOMVJjKpXYxVg7ZGRECUKDgTcuFwJ
xpMKMVbR3reaACEA7HBZDYWgkC+BjxPWw7HVyHETjVtnOeUIqDnpJ3UMJnsivXS87Hvbdq4MtHLF
wv32Qz+1fbulKXnObvUhn43GG+dSypGpqxhet2zn+n0Fdodce3QD12TMgMc0vS3EYJrcXRw/j99k
nFNADddikaqtNIZbrIF1noU0QZGKzjYaFfnDLRQ3vqkrSML5F/+uzIC90GgOLTKvDdsLOntq2CSw
inuyUNziez9w8nesIGOym6NZMhUTXHUtNjRN2jw4ZRcJv0turV2vxeIjJ7fZuu2Any1WCwdz4eBt
NgNzyi4gmEb++rxwRrRm27+cUEeOwQYSSYxHO4dFs97tHq0NpDaEGm71epgNR99PmGwr1Fjdcm1Y
8ky3okIpxrILmdEN+WU95YKM7JTlUNNCFeIhaUXIkioLdeH3eJ37mpeHKzwm37duXOL3zkv6F36J
g9LjHmZHn/z9nU+5sVFdNIXNnWXCzUVFvZJnqN457DFHfX7vy4pZisErpih5fndnNb+5k0UxSnAg
54CfhlHI1isGS5x7E3kGNGLQq4lNcXjbQdRVknJGvoBdMFU1bgo77zKVIZoFiiuXrPaKoq9xwf5d
kTP9Nt4oSBG0lgNy9HpQ073EU3h79rH2cs87QaWwTIkIeotHhGzZDCQlMfotMB1mRTvHYCoPSu4w
fpRELNLbr57iBnbTByFGRn2ReIKrhNntkbUQB6S3QGbYQEOes9NGiz1GWg0Vgua0gbmeWgdUt3A/
so6J6XK1PlJyOF6HCsm63kfPTZp9Afk8o4Ke3QAfoNBiXrXCEbIcCGm2KVqabbn55O5JR3Qf3wgC
N3Xhx8gdRQBHR6aggf/Q79HIKhuzL2gVyYN2dbpX0Hv2TF3IiSmYHNeDaso0+dF4bOmSQuhQSR2n
mh0Iy3qtJeCVnmv7vAecLZ7ryPtGoADFvJpuKQGyN5XBfrpsgfDKjOl40vKSFyEq1PpAXsZDfLhe
B+fLGZCRbazkE6lw7xA7TsbJNBoe/4WWOSDsLmJVEFqrBG7c6i9a8SdgemdTbwGyxOMlDhW1zmwa
2MG48SbTOtXS/QtPGyf37NyKWPjpsi6kLodx5cJh8xZJAgsilO+4ct/I7UR45I06D/OtnhGO5gOG
RIDW6iSCUGAfbUAdYvQnS99hJjo++iQC/f0vTRZWZOX8VHn7kGKc2OZJbx06kFzi9X5Hm1fFYVRr
6dq7xoeb1lxFs3iqONBw8QtMfg51RvkK/+YwuFbysVmFI+VyNIET2tm9ILRjQjq4wha6hlpC46wr
QVf5snF9QZjSGCVIqRnZf72c/7m1pwpFE2XpJGiEZPPRofeGLk/QBSCsczQ1Q8qowHpHBn6udLX2
V0lbgVv7ZcU649Vi2N4tpXHaId9ZMWETtTslHQD1r28Wo4bOpywiSYj1/GzmpbwUfj/r+T0sRXfB
KWhSmP0ZuOJ6fpxYIGVWGs/sCdV1mPZhPmLyatIL0KeRuu7XbsTAE128p6QjFqDfUrAdGQz+DB+m
PFdkAgWZw7s3bTUGZcyDcN/OW6xK5/U0OjvjznIh6ZArw4LIJGnncwLZZW764KH1SJDXO3udLJvi
CRSA+xdI7ZiHjLdgGH4RnQGx5bttMdgl05WPtnJ2top+WaZqA7xlYU2TFAClwvmLcbBchRCWvGNS
49w+T3/E+Vk+lLo4mHP7vArA4SDL8rSLCJq0bmYmU6aPkLMdQytRQi6phoim6G+OAvI5lge8xn/T
IVA6gZOSkhhJU4eCcBI2rj3i0MZiP0SXQ6bbE96ihZR8RQl2ACQU/hj4NizXdjUsv2r41MOdRexS
kHZygOwYIPaSZvSedWiceTsyLQReayXAr2RuKBMXyaPBca2T/aEz5zlRp2BF8kNorTEfoHH0vBOH
DeytG+k8s0siTqg/aD5RG1GUn+JarBtAOHSqx1/aI3x51x/WG30nBnmmnI8S+ZUgp43u8tRqIQDn
JHZXVu0bkGKAYoUU+OIk6BHVXcIYKwoYex8qIu5DVkapKX2ESMXnyTOI3T6CHhsoaiM/vETbkYUc
q0xGiVheUC34yF5DWpCPFrNoQAuvrfag5P5SNTLxXFTQewKbZzR8LUsDij8tBCA6DQQVRyxYiuqp
QzD8tb+FYjz1K/7irEe4tGO+VNcY9wqpmtbOsuY3wFQWevxypQKFYVWs+rAym85GIN2eqN93EYZH
sRHG1dv33LIJvz8EZ3cPGttEFQz2Z6yyFmc28Zg6Zwud5ZvehPnTzP8CUbSIpI+U7KHajwvACyQd
9ZpSBzqtePkStXNhTfrBn7OGmX5zRbwnk0i38TrvhiAZPMparWWBVNXQ4VASp4f11bpVEaWc4qMw
vPhRXcKnqW6mqPnqEi+isK3bXQnhj5/iV1w4aTgiFsqYPQoSOncm+zjU0i1GHnEtGSO66C3jLgol
tAE6t5WuhoFCzILCPBUradR29Hh5BwOFAUWyAAHiuVfIcGVqXxK0NWAybsBr5qmj+32K8VtakHAk
87r17mOKW9XkMMhZ1J5OAmOvjtLD6fC/Efa7SnKcGlW6euTDbPRj2/1TSs3dOVZIMfT24Y+SQNl4
Y3g2qdjVNydUT6pVBZl8NeCzUIof39Eqc0tCBGYGzzrNGjt1CRcl3Pcy5LAW4ia3jI3nDysUEnQV
m4UFjbuMQcj4Lp8pznEj3MPr1/bxLIiuKbyJJ2detOdQhZ1i2uN1TaMQpJXs6Ci0Sm3T/M5wH5PB
eqhlSPjGxpJ8y8HVBbj80541n3PwhZOnSi6i7Pq8kTFdPTij6UfqGRO4Dy/YlZwui8CzNA6zfb85
KDdc36bhWKR9jCUfBexIU/sz1bvolgPowPn0ehwrnE+r+nBV08aOYIi6qSjokET3CcFeiA9YXJ1F
rBCr2JMmWj/3UEVqkOKL3vL+lze6m7ozKqFmtDOABI1No65SMwenxwd/axwdS6D6AgYNCzdmqkqC
e3yNTnmDZ13G+0EYR+cNn7K5F/oVQoKB/gSDQAdDtkES+An/gKzIYy+zxvF2ms+N4CdE5g7xW/T9
1WdzM+kNqLgfqWjhCbvcBReTSuBFw+sdTlvAWU6kClYenEXFsFBJHihrHcDwMnx0QFp1C4pKamHT
BUAXgzRGqtLou2gUOxBBfzbqw6BRsvvpu7YO+AkfbSgbAOLAiz2oPU6IhXCAXdv0SS/2avYX5iA5
h8jmPSS1fEdti65MZDtC4hnevvabyPTie+yNnZh/0hlhdY6hz1PVa0u+i7rzrZhlETlQlpTAH/EW
GR1srzslzr4iNpoyH7fpwudmY3Ofz7TgHMu12stb+9BK5OStjrIap7zJp+2NREBbz68Yh3MvDGYw
OSwySe0ztukgdoYe/mwZZ3DIWyn6OoAoCZlyHzW0/+BhuyXONZBfiTLP15x86Sej3D/c2QEu++wO
5gezjCKp8OhT7mqpeHh6tx18riZ4jc4qMbNRaQMlr1PHn/QtE00o+EErO735G23t01bTKPmnFJvo
Vd1/YMxzJLPw/A9mnxlPVXXEaXtgVD6McJ9ya9XD2WcDj33caYuVhsGu7+sxzIaeY2gt+NzTkvKT
/MgjzOB82HhVnHTQlEuEWHgEtWJN/6pyA6MU8AjFDbla9AivW8z6vkWSVzUuVRRJ7+LtWx+3a5GE
Z6rjY3zBpKId3bnDaiwzQYjygbhn93gJfCR2T5sWpgbjV5J8yNzJ09qMoEGRcMbEuXMm6i6Hb5YY
WJ/pjPbGhAl0yrr1XwHQpjk5tfkGKQzmV+EUmxKM9ojHnLRI5u6yT/ohz84wuWvFkqlsjmx8ZsAP
xmpg/O4f/IEbOPYmsU9jCB3sMWxEmCdChQlgBMAlr7FvOnDFje02SvlO57zkIugoteYaJ9OSq6pK
QvlpoBuBksVnRUQdYfrYgl8VoUQ1r8ZJq5BgjDu4cPDmKON1AkbHtG4eAkMOJ3fUcgIdPc349Fcv
KxJlBPJRf4aOvXvmAJmnS48/ydJo/H4Q7USyNNnyzapZjxnBFj8HTp0ZD0qK4xDlbpvymyrx8dM9
mQHraXKSn5SsUeJ9NaMNEmOpCxLLG3KzB8sKcxD+wIi6cocpy6xVp0sL+qQwy2WZUlUNVCf1534M
GSGoLjJawdVy7dnlCdQ05ck4aNEv2ecrvWg1ayzQ8iRktX1GNKuk6WTlVwgV736f0jY4CpR0WdVZ
AEIFj+lojly+APD23oChpqAtcBd8KIuLW+uiHMCxwYafPSgcQpF4Wf+YR1qHweScbDbP1DzuU5Jk
E5uOHgDzJ4canbNn1QglL2HM3HwY2/k58l/ZB8xWUco9L5HqoVhQtFm+Jmtol+iEOqQ2d0cag/2e
1OMWk0n8a5EFOzTKIpZwvqObE7DveSzk3d7viMn9I2tF5ogeotUh1SZoboPJ+C+4hG2jWDNMaxEB
wYzbXQA5TIRJAzuhK+lCb+O368RK3GPjO8xb7vH1y0yHbEQcfzczaiySSKM69UivPjwaSspUbgRD
82KGN9KkAVuG9ECBUbSgXaPlCaslcxgEp5CQpMVxoUPCTn55rqCXZh/CRmEAxXE+P1QlOxYjRZ46
tFcDb0WAbxWgJ3oxKy7rpy5fKAFDQzdhy58W5/ff4SwK9FX+cM2jUMR0jAkaKfE4FLghXcGrxQG1
JQzpJvIhmhwsY0dnbcYIuZJaOfvz5NI+lpfGeJNE2sL8hFemObFD4psF48lZY7A63QEZpWonGsDp
WMu7vXb/jHKRPhWzwvVYeKE507RPj1Lm+TKRjtbxVx4Ez+fNud+Xrn+Rdp70Je5zsA6qFKxuzDnZ
mWOr3LTUkBxM0Bsl+wybTa/DrmwuTfSVM/ylV/JbKZ88GztdUzc+ZLpWBoFkvlYlWekTBD59rfRJ
x7SCa542V8PNoS1l4jit8MqHSncZYYjpgQqdzZ1tARLl0lzzKGeguXuCAeMm1m2LTCONH1XHIQbm
BYMlqKbwmn5nj5HB/JQdVF9NdHqv1yUwSjMnX6HizWOH5qRlXto0ibsXuLqWvBzhetT5VzvCh8Sd
zTI0YsJbX9AF8UJECSKNDVxDUAkZiMQpEPVKJwl8NZVThr4hZCPCoJAj8nHiDKgFp/uLNNWlZjh1
ELKdYox74SWKoVIBERv047Z/mRPLXuaKxf3UaEyZau3QOabdxVy8mzG6TlIOmGas4ZHw8k+tTa+Y
GpOiH3khDYXmPeLJdMZ+PMV3sohKD1GuL5RDZOIc4NS7iSGmAcwvQ+gg8NaYFztprobJhKzc2LzL
juh+HjiaAu5u4EebKlwkt0g+W4sOPiF4uLxq5ydBt+UQZcdFxpvUWheJO1UZuC7/V9rnBHslGbM9
5AgU8GyETx1pVbD4xuDZBgwo4g+9R6/ba7vc4IT0F/TtsZO2tzOoogAiMlsZnZoi7A6Gbw765bsY
4pCTV+ifdKrTBXCrKA84ytrejzdTnPZcf1jXDOTRPBWZzB+spNOE0b21JnE9DXSkXeV+zGpf7hzE
ashMUFbh5ZM4wcjrmERiRotJHyagB4n2DWBQDnAfvHvGTmaLCci6smF2E1mA3TpqRXNGzEVu20Bz
2+HGQjRlAsgoAvcgnVeSjVFsUMpLnxtWkczvqUeGtaSJn24eRwujsdaS5nEi28ShZBi4ELrzmfwM
Ph86XjE1gKGkR+JiW2PDLl7kusvMj6kHBdPmSVmAlR/8t0PtNr7Jso/J4bSv+3nc89plbZaVPjnr
v23zZYBk2tBA0jhdKtjuXLurl4LCZrrCFOlo00W/hpXMbWNnlHhIEF9Vcj/bRWjfh6+Uav5S2Ied
os8oVN1hAi/tY5ea3ki0Nte0OSx+kFYY6MvoIzOHunBtODkPravo2ZnoDDKXAkCKwYHT1/3gUVVg
+0JJoBYMvXg0f/LK7+05gdcdwZbt8/EDi6PMYvamhp+8eIjfG43De12TIxWWjrNUxqmKXg6lyjPC
OFbKaKJFgf+Kud6NSvDOwh5Bf+z4EttiXsnUn9VQvh6qf45fWxTtF26SbLIUtjDGR3fO1/xYAQgn
egZ1Z70XeMclNwIAO1/ghAlAcQOqdw3irGmCsELTwi8nEKwXGgCYVWlv70s0oALqiPRPTgxs1vt8
9dtYKkewff1HLOJ6EQIDNIzCjFIVb3IZvweRG5keE70qDGMpzsygQOhMSN5IBRkeQeduemzDYNoI
C4apQZZAnGo+9/sVt9vq67RyM9X3K8trk0LyGOpz0SQFl9e0VIXOV+DcHiD3+36vswhHJ+7JPsQR
wwuJtgy8Gexw2nthaLeeMvoDSXfHeujp6ilBRFnL/OkmwlABkLLSKj1r2n0m0KjkNQwt6rMnRvFX
WKHC2JjFfcZZ/MZTcRuxwxeovNpYcrM17gKQNFKeWdvplJZBCxu0LHKO4qW8qVt7cuyAOTaF3qA6
xEptnceTXtjt+5v4UI5ySkfHdVUl0XwNcB+KVrEuGkJ+SXZy7yPD1t5QItA2cq0Pb/JTLnQPemd+
2YOZkY438hYT81RRFon06SB+uSz93QDGo0fE/PjeQUkfBnwY7UOqz+sDxgr8DWpCICdHGAHynElc
0zDfupEeehRz4oyME9MxYlHw805K+fvOrppPqmEviejIFx4blK3FVWZnnWNmOubWh1CYW4acV+c2
lcc+OdIgyI5fsrS9Gu56h8hukoR6NQtE7L7S+4ZOCSw3KdmXg0jSZv7H/bnMGDs1VrTDTP+Qsnor
/3av1svhvVH5NW4yoiqCnmv/Tk+w7wmoDvKIGxft3JCvTU/dwORSBbzn5KZcafAjEvG2NPWYPkbv
QmIhxFQWBnycqT4Cr+mGbphHlAv1ZO9/mBK/DuIDLUNgw2jEBIRRNXs9ZAlBAhIpeA6YPhpon7Q2
di4MtEesLv75A9GsEFyAD/CnNjFxYHS3KYVePhXgFN+gfhaKTvklfqrp4lbs+CkJFF4s7EdmplXZ
eefqLqV6C6+Aak3rY3JwfGj4GC1inBnHNZNS/bI3c9nvjRR0sDw7Kobh0F/YSb+AV94OlEl1x/V3
ShUcicZD98EcIBqc0NLJb40FEcv5UtPMBX+9W7VheB/9YVTGAGsbIJSI9Osq53zJ2Tyk6cD73P5l
3gIVZWRqnrw/O8/DHo8acH3+2vPvlHAqlaxYxb8JWXuaf7bc/q8cSCf16vlJdnR+OLY63Jt7iHLn
oDR1N8n0F91OQmp1dEnDvMXjPN7VnW6sl4ceuRuTd0KHpg0M/RmIyMASxUBJYRlCQF0VZ5wKFEdo
e3yTmM1f7cjaH8Sky3ZR0vn61mjWgFgzOdUcMdOEwueBkxty9OQa/aKhXG6Y1KZl2PmJaYSlaTwH
5aOBQS4rdBwaJORkXGMfCMiZalqUl1RWUepcH9uCAA2GvnOgXM8fkx6LMl9/QB3sowrqSXhaQh80
QIvcufr3WI3BLIDrb2BBnMMO7gTWcQ+KcNp4o/TSqkqKn47wodqCp7opm9gkWIXw/6UV7d5FZm33
dVXEH8vbt1h03Kv0PyEd4d31EhKjiC3f8SjyAzE7YEq+T+0Ki4B5SXqBz19uvRt6DjUg7v0cqZMW
otI+ZvH69aFFwiH9ynS165QB8B37Z/+3rKhQaSR818sDeC5CBjeLikCSWZwtIO00RlVH6jpi5hnn
LkHT1Kwhkfj3Joqhq/Exli3iOzH9s4WVPQHsbq8bEDuJRDJgy8cU6SQSTEGkqO7Okp/znAmudc1F
ODwLFsTtyX8rCElGvcED1Hsb+bycE7QmXmzeRpkvtF4Ms67u14iUNjkZjTfqkIu5Yi081zb7kKrm
DlXgy3uL+isRNZG4R47NKtqkQ2Zuv6TKRo/pNr3yv/drLW26JhB/RgpaUIGF4aFPT6gfQ+Qap4QC
USnPCZYr0yEepO7dlJWlTTlbvD3wKoaZzwPtjae86/hMPN13Kcjty/WUqU/q6i8S+ymdlJgfZ+7d
Kae5AukxqUmsGOpvnCda/JfLWtJqCIWysKKiu5cfoeQ1NWIVdIWPEfyyz0jOrUFZEgHKCj4aXFOj
dlhm2HHmGAJit9RBZm5LNGenXvYwibci4DZtTG2pgAlginbVRL5D9Bkp7efP2A7LJcaNB2CI7kcO
binVd6QcbKebIFrRG3iF6iSlDN63l/+9aGaghQgSiPwXRzHixa8Fl3Nb+Iel4LijzgaNuXVSF6yS
ew4CZiQoesrMlxm2+gDT1LLBB1BHyEpiBqXBK9E010zpst2D8M6LejQetumftJVaOkqQMA5+oaFQ
ISkQvIPaKJw69jmJxStbXTI2HugcAc96xWzVywaO8L+yn2T83X2rKS4W6q3AL16PezvvAAsBjNLA
lCTI/uKqb/Q2O/wevHPT0pWx2s2MW9CLcCdXajBJzO+ghtneNI+HWV9ecLcKZk3wrYfABCW1hXVx
ejqSnO89Jj1JgtdcffWN4RSVx5od7oCvKegUkFTZ0zTo6yp8PKp0Am1n+QYvDO5Bfl5rc13F/ZS1
SmUo/ymwONjTVWALEUhQONAm0K8IXThgBTS2Cmp9C7jDfDH8LABU3o62LZwfha6kut/6CvOfxG69
ZznrB2PdAU7G1iP1GeOYta1YzTyO9Ey2b97DUMUuL2hkYsvYhI+a+pTZIhBDQwcY+OEOD/8aEhj6
VobfJot4YnMuMqfYJKDLFHdWuW3yRTmW1zGK2uFdHcsXdwEFppvjfgKGWAbV/XzK+ut+ubugC/k6
jRQEqJtosXfJeQy0Tiiwtcax3T2ZgBxJwCAKwB426uR4RVF0U3np/90nwZ54EdXdDGB7dr2mvxc2
jLWjenzK9E0ilG6tA4iAjw+V4hMYoHGvZq1BAokPS0WEQKBtYI8CaHG862eR04P6GMj6JG2USw9s
OAechxHVz4iYfy3bMQFkmyx5TadRAZxuYlLc/Ei7Swupeu210hnaZAc81turiZ57EyPbQo9bvBCd
UvzejwUE59beGtZ/IUsPPttaiZl2o+qagE4tXeDzP5MonLfU38T7TWg6QGx8lCIbVrysLfMToVOc
N73xIW+tJpIXggjif9bTNg3oaDHOKvFDqyae2RHuUyv0RvnINlE89I8UeL6AH7S0p0BOnEoslUUC
EXw2bmp1SyjvSsfCvwq3rckK0UBuWttGt8i6fB4963jZIC2D4kJnQSnNImfSAItRQLjzxjYWWusE
bv7JP21d8v+wIwTHStrjLx7GhjV5ooHOKiyLqSYiVXieGtZ0V6eOeLCXbXLd70XThzuK43QlLH3I
WsbfSdnjRdlX8hlsvsljhj19vub59wq0qbG5FOZRIEVOJStMmD36V3m1ZUWZQoun1O3SZ8J3E94q
E8JWH5ubfA1eSX02KFKGwqxHOOkebFwjmFSFiMWI9AZumBSnnJQ55vLw9VHnrwsK1TPvz4Bl4D67
U2XmoeTnc+aGXrWuKg5M8Sq5sxkMbc+/CYUDCaLw0K2Al4YzDCt3Og6X4d544yhd3d8fAfnoY4tm
BSB+75P2JwpR7c6T0OCjE47fRJ6hWCcJgdOcbaytd6JMGuxHwCQO+J8fuEQmPf0zbCC3weTEgUzK
Dh9skMqSlCCYtD9yKoSex8G15jJS/HeqvijKc4LG4JN/nJI7cFiq1zAfG7Q9xkmVz91F54CwThvS
JIHmRcx+0sUsHH6bi5KGLbjTdbDn1gTYgLZpJc0YhbmbCVjoDmTdca8gn3zaPjt2YtS0+7Z2Yo6E
cbxyXloZUX3jTH6HMfA1oJ5NMSnk4WnvYFmUhzqxtpmBELMJ80Rj+6ZfGNm/WXeKnELFfKeZP2f8
vhLDBprBqufa2VSAJw+kD+xFgtf5hI+kSUfgfwsYyAC5ajR1YXdfQkBT0oWAyyhPYtVGmS0dsrus
mbC6udt+KXBSnJF54+O/TnAOHZljNX0uXsYF2g/Qst/A3eLLQk9mspkzMkO2aBVb97XaS+BMLvRt
my4wmUgLQcTpCsylZSj44mMQan8xn/JziNlGmTHffgRKRSg3fzq9gTQhjbRWr3ULe0LSbUaIE4rR
yL4CbUPNFC8hAhesjWRgYDf304tkbNrtiA8qrpeHP8mN4Q2OmvxrWBrTmtwQ1wZHV5skkS6/epQq
CNJdfXqB/xO8qoQE4q5vhcexlJSkN/LPjT2nx/m5VZzv1AUDhrGRD99ld1HB39a/RyL0ye6b8e35
2gu36MgeTZPz1bdE33LfQLP/8GUT8o7di0ucRbeOyHdPk5Kt4tB+ffArOtSgvWgP8AmyOGhHvyv4
XC3ZQUEoqPY8MUm050Jk+GAgmJDDwTvAn/ST6YlIsplhPPKZ3uRzJatpOicP4i0o+iSxKTeETKZF
doojCwYlBSB3STYED1j0mf2CbbH1JC/Zl1y3h7fZtE0TcByDGvQ+qWtw4N9kzne47ywlhDENGT1k
q2Dds6P15bS0tt/U3ngb9Y/re6Uc34VS7H0TH4LPOsAgPMvPdHmF84GiUKT+uTMU9wT3PNjFJ+1o
u3LqKANotxzkYCeJ655A+tm7p8+O6mOtkgZ1TkO8PU921CnKPmhHxobtF7u+385OaegmRD4weBQn
3RtQ7Y65ARvBK2YcvlDGmQ2L+0qi6I7ztlG2ynyqLYuPezEFNMQzKF72A0BPYfBvtvqMJmpYinA6
8BKApWOy7z44vT1c1a27X/SJjbkfTPdICYgIVWc15fPKXH78CytfNMXCHipE8pep0015jM6YbyZU
KVXwniRBtjnUS/Blg/TkeUMkBYjpp/+NOmdNV6P13JDhShbvLr06N9LE/6/gRoV5vJ6BbMpyog+N
hFIlu7r1U45aIeizf+655KgKKvSW67nbVofYOvMJqLFWVy6+q/pSGaUuIO29YTDvOx3Rgjf/7dZT
OZPEyzoFG6hq8HAjBLclwSjQelUh/WvQDAWAmpjXn4o9VSbqyM+0dBYl/tO7X8e5X8rTq98+JkgP
PgUHD8Rdvyvj1EINxuX5V/de3BH2JC1RVLvDpSlVrbxUju/+th2y8jtSBxuq/1qUh38KsUBjRyKE
7TgcQcWVvW6ZyWK6ia7UUWmXV9hcEzCCBcZEDB6216F9DbN+/ykiTaq8Lsh6qXLu+AT5vajCt8zj
ovLUbWFvNd+LflA6JeM7cerY/5Vx8+rhjtsAaD8t7vA6Df7l8DHKf93fWYv514GjZyUamgM8uGxW
0HPQvK1KaTbGi7koOMPa/iWTxP6oBUX4jPY9vIF21p7M/GzdcH658u8Hkv17+aAtheaRVybmH9jK
YQKyGdwjL95YAthYak5Qs/2/jnaiTCsiuq6keE8wXpUc+Qo2I9K60SU5H6LfNnuf7dg5/IziP98y
lLyit+39ntnt7ow1N1bDnkeJEDW7cWP5rDx1hMqy7Zs5oX2A7inqf1IphbGcJsCm17w13g9e0ccF
aaQ5aEGFSUkeYrDWfGN8xB/iYsUcAUBqalo9xrWZbOz6mgKLMsbxJ1V25ngsp524zMRIMO+IkNEu
rDvPmpJwCDo0A/yXsHZs1Oyr4HmNY+tRsprp1hHSucJr1DvZ5NaNP/1x8crLDgeld6du2NoSh/p2
geAKtFCDQXz4kFBrF/vVf48sM5ZAfinOs2U5EtJX6th3jf1qpYQgSc2JfW4yS7H241XTlUQTfQic
L1AKkRoGOgEFnX7jHI/f+fn9g6VnjmbOFueLRQa02GqXQzi35HgFOm7K8NEzDKMVFsBZxtef1SFB
9UBWbRw+iCdqFyoBXWLKrhhcg/6ydmnWf/QDloMdn5lv3a4yl5HpMEQTVmBg32n5MQgtkr5FF0Sr
9tr3I69nWLc+Sw2CnJtGUp/NiAAL43Y82AFKMIfHruhcRtRiYVDLSYJUvEc6cf4q7TncT1mc/20U
YPoHqO8VMlGh5uXOLjlrvPTeE4L7cYUzi9bY7wwZkJFOpVdihDkSTelMxXiCLNAR+FOJE98c1qMh
kzR2trNjuuVQxyyeDsNVjXX/7R7vBDA6GW+tfK1WXsabA5Mf+6LWXCeYEcAW22p4NCmhplztDn5q
VoOXtWMz8hd0KHHK++XhF1WusyGh95Y123TCr804+VLTJoKujRSUu02UjUA4AG4ejtQxwwlpv6sK
d1wacWWcnBsVd0bzqDbSJIVyRLF8qbEB0MWBmZTornwoxRfRDZtl1yZ4yheMED1hWIkjqjkavS3H
RkACWNMdUT3lUEMuDJ88GOF5aHVWSEcFFZKrAc7dXwJCwMigx9ja0+aszf2bO8ebubDsjdz7e4bm
j6wl+GFIxIsedydVRSO57VZ8NfYJM5P4i/+x5xCKVA6kowMN+irKnNYzKEcADej8nnHM8sFAvhZe
Xq8gy/+kEMI0EnwqFyUg8p4vl6aG7+gRkt6JsDpN5n83TrlaUQw4uNLE9ttJbWci/v8ID/r5PUYD
nJ4g+J/zDQe7Xln2mRxgz26fogtPlQaUaIzaeoN4M8TG8Mqe4c3OFpsY3GUyYam0q6Y1m1VaV8il
atGgOASKFVGVaJh43YJdQUzRqII3PKyNkUBxObyb9Gx6VYE1RCfbM78bioKXuiXkGfQ0rUOMYRwm
TNYROTbF+c82ppVMdXJJpYMfaWdjogwtB1L/nmYZr465obwjz9U2cNDfFr7y03rqkrXka8otBb5x
eTqyrXk+Y0NsTl1eRQlzkNgc60NMXZyoBcJzj3FqfAzXX/+W2qO1E2/JwqZhdo0rHY1MG3+spU2Z
oG5NEeRlSRFZnqEwzVLGkffQdCJLD6x3XyPqzXU0tZGcM0Vq92LXv/+hCbdyVIL9WX9hF2CaO547
n5Yn9N9Aq7W76EBC26MkRIP9RqnWMYEjTByo65CnWvsurMLRIhxa59/ZRH7nLrzsRXMjSym++Uie
5ro1rneJ3NuFy1WgVekCSq5+Lk34gBe+YcN0pdjlbvRqoZZK9Agk0jcRgpMq3boRak6F7PxU2iHV
PJPBy146T1awbbwiFH3oGFAr4v3GqXD3YJExas9sIYvfR6zLazYO6gW0Y7Z5il8AkHaulDVylP3E
aZ9o6jsARSUY6Ir6UQo/r3HxqJnJDPhJgOnJxtES9wtdGxevvPpAOOF9BuJeDDRANvncWRVxXilA
mZo/3illc3iZgxyl9UDSiYXjfZoJl/1BpxpbygtAUu76N+ads3IoNgEuTl8XI5MZcJFagIyTVLPv
P87vlEMqNrtM3jOleHM8PKUX+JHtH7+gm3ZE1+ITyANOd6N5jjgihyfVGHD02znW5faRSxgaqwRh
8ccrFGIwXtoLyH4T8qOu15H16SPEmAwLoNHmPI+KeVsrLIA03BgqW9BggCgW4X5HVpIXFZRGAVmb
yGvkIgxC1gFoo2WmTyyKMN1uBRfa5ISLB00giqNMx6D6TP1p8sLu7TPIixYzy74jKJLQ2zeCD5A8
jQFlAPAE66kG1FQ2qzl3ozuWeiiVMxT/LyCwgV/TvfrxdzGuSb9RDat/Mjo3d0cOkZZPqfzOBjh5
IHabL8j+zx8uDABtRBSKbkT5LOz0xJV9D8vGSeCtVU6GWLXGsHXl1hdQ24THPQJibpojt9jnWkKv
eYRHE+2a0TPqyE0KWsP7fgMB5OSbxNXcnNLcEOwFT9NfAWzIa4HPJRTYIcrkJsu35edIwmpYl0eA
EA0/S9OZ5bW7ODyJ+9e6CrMah6MH2Dpfwd4SAXv3n4HHs9b/HD90n/gmO5qu9Islng6hII1OdojW
AcolhWeXymKSoCS9KeqpSBLDOGT6gGLQG/KV3nwrN0xAubkXJnEUbZeveE4wfAFDwH06OgHhIPQP
+mDzQ+jvrB2DXblh9mhKkK9k9ag92atTqxeVLX2He+m0jnYtjveaKC0iC09CDfeDIJVe/BvJZ10m
PpZWlgooKmGcPwMXtcwz5MRVvfmKrkJa4iOYVFj8VIHKL/UNpjpF2pcy5ceLlaykzvry1KJH/SRw
zm5TpWJ2anmC9/jhA2lWHnYbeZ3cXsH2fLOBsu8RkQC11Bw/t2rl/dMXrg4Du081jBiRagnnA0gQ
f20oRqQG8zOi7r+pI+rAUzV2b7yR6hja/YuN0sP/ksp0JYFXl3n731njoWHDPKrwx4qxuP8MIcru
2qNzdn9wu+kIuFfwR/5L8C0q4MFgilIt11/zRpoD57ft6cqUUEB/xpwizY5zKzssF88WWnZmkEgR
2Xjp6kgdasn5qvvaUDzs1y+xarjy/1pa7Zbt5iFZXFJEPp+dLQKHWU5Hu+P/MCgVVu2uEa9VHYm8
ded8d1EynsTVt92oUh5qPTOgA5sliCcTAk5vSGeDkvrpWkw1hHS+7514r589lRuY+M1eSbBQz5R5
xNlj6Vfimi6ikqRk5kIiYsQYcruqn/SAEgKUZYPtFz6TlNV9eOuG45jr9gGjvHy+3c9TBNL8jZUr
uCbW1E/k60jc9g3xNrB0dVCzOz474lqnZQZ+UVRRP6+dyZywl8ciksjN/Y4AyWuFXt5Z6nGCZ5bo
fk1V7l9GPRf830DtgzlTPqjuav3nLX7F+EvEh1d2Lu7SFfkxpyABBEXCR/fvISd9a4gS5mWzEOaQ
UumAwgqgMVde3z76PgYVwroexzH9oqkkB0oW2B/nhabe+IOnVohS4RA5hxQSuVgi8uSO2FUTnaYL
opHs1dSleMidY2/HMF61h+6GdEVTeqBWNexuscHS4umSR6S8IiA8Y2IoMpMZXi6S43SbJCm70K6E
vhMBOyvWbOgX1lvyVD2dn67XBN4p08U/ybpl4neCrLRoCZ+RLd63l1rVn84qFO9SYuFZdHYbWv2k
nhQdevMK9eqKF/u8KJi51fJ+htwdkjUTheOv3/dOwuNnd4CtWSkSrU1nV8Ugwmjd/Gw5S69nbyA6
oknf0+gyJMWE4BAQs+Jfi9IOzoN6tnEIStXT1SZnG/o5nEI06x4e+tm4CRxEdJNLoD1XhZfdc0hp
zXPmn3vrsRjYCYKkaA+cD1qjyFi4k1h79KtxmfhoDwDIeuX7GrqQRJh74y7MpXpbI6TAFdlBvhrR
7mnoIDp3tP5Zz1+nSjZ42LQ7S4LYZh5Mep2VSyxb76rKz37GwCgozIMuXThsmQeCwd22DHPKkkRB
xvgNzChWTgV3Aaq5fe8HJzosInnMz1Uv5rKP+ACtXX3ajzcMR/LBsLIL56V8uQ7AG6UAtq892GnE
CZ4ctGNY+kF+qkikMoDdeN/BGgI53sk+tx2qzxRQo50lJtMjnWZejy332vgRJ3c2CvD229InAZDv
26W2D9zZZO7rTJ+sw5hOO57WhRulAgkZ/YgHPoatVpnX/kd0R5itShal6GNZ8ZmoLchpFU8e1/n/
7azJlv7mqt5TMKWjA5z08nSrNXx1C0YSToXooEJQIxk6V0gtFR3b94L7ZpPQe4ypB5tuTAhCMk5t
aStfNyu85em6xQvoeA7/IOdJ/QoTOXPafu/VFNy4xneEf5RIilNqNJqABWnruOg7SzHmIeW+jf+t
3mQj8mXc/ipZ5uCV62wScQ3VgH1dGIiZ+yKTlnE0KjUtgpMRfekfNgP680M+PrWzzK2o+pLLAf9o
6YFrvfXCLlBse6avXGoFqfR4bPlv54N5aSw0e3a4ASO/ENC3D0UormiyfmoVWLvY/6lJWiVMKE9z
b6ifrGzSEZX5v9jO4b8lXsJg25ZO1KFFnBNQLS09gEDpF8TI+50esVugalxtYYrszUPxpyUyMSZJ
MUH66FKX2fjbgJtZZ6KvE53fV5r2eTKBmxlnood9h3mC8tr4W0FPXHnxNjj3jLzqekNrtQKVkds0
kanEeAf66Rxli6/xPEPsG+ydA+lzNf6xs9fSiPhShxBAYfJeTvhKWfmyjZ37gGyZv1eg8JpCVskl
tyuSKhF/yD4T5tqphVZUMNQd2OK7y7zSgHcEqBweYMzOHEePbSohkysqM5Uhst9gGy4sfZshliXT
JuDAVrE91xD4Ga/QJLapacVGsZTc23XR11EkcDu3F56MeQ3oWyDATmpB8IrwVmNHB8EzFMglClU4
w/8sSeY+lCc5vSOQbjIR4ah7tR5Kt5ZIvDbTQOnreMYRzZjDj+nZ+kFBsETxIypz0NYi+4flzoCb
sO3G8sFBuQtNSiimElWk6KLauALXxQstAhE66syo+iFEvisaNyupCOJ71eK9wISDuRrc1sgG7+I5
lAeVqALlfMx0JFIkesMmrtOdB4ZL9HbuP8fWMAlzX+v9bHuFy7y3HWjHCoD+uO3rwAcRU7SMoD/u
6M0T4S6Ey32O1E0BFvIbfaKmpk9POnWPio6R1elhkSf4KFvWNLwiL7rv04rilCJmmrnk+TnJu37a
auGzDCzN1HuamMr3U5ogZVv+xF6z1fer6wfAvzV9a9/u+fGQTFtolwj6dgXcFzBCrM5fBJH8+fiX
JwqQUdgf81dlPDJLqDtq/MAq9sIDHhX3F2a/UBycAQQZ6olykaN/lKsLn4HEu0ZuUAseYr90FXvw
8O17MAU8xhS5IhMhJ+sZA/6UVGLat6UxCUFbbpw7cnyCF/TGqqDKJhZ/AZW818816Jb0nk3Vwmm3
KoVdN3+iGUsgSHGUFrclubtZ2V57fZTKA8BR48oSgPqviM52CceRUtae0UVnpXdb/s//auMdhOzW
TIYLyhOcUalO7B0+NcosUDN+Z5znFT0vXndmdjfBi+nRX2qlmbbsv/BQfvYbaZk4vi8dcHlSlRxT
/Kx2W0qCdBNri7Rr2e7p31Q7OO13lFp5SwzEdZpo8heGYREOiff9zzQXA+hwt05XFSp4fTR+a3nv
3gKTXtbwpG1hl2D+HzCmvYPknXGj9LL04635W4v/exNFv/xvTBtr+wxCAPuTBDGixom6Dz6FfMOo
eSQHHcQmlB1XbQH/vfvfaWVNzFfSbNZbKNpvL2ye5Sv04K3LY+sZ3Zd5qfca3KJd06m1EXoDRhud
D0G0OUshzZN+1mQyr3M1cov6+FRDzvLcy0jHqIkoAGauuLbyrLF4cNwRBqnW4GnwXqdmhNAKtXCG
rfMM9uctkQBkmqG7CuS1HhVSDAQaSs1Jj3bnD0eCe4QEcZTjwU5NsJvbFr9I/otwA8P1IXWhKBSb
ENCge4Qxf3pgVbqTiUkk/8v83oiyyzxi6N2uxz6pbDawQsvVoFTZ/mDvZRypRTdtGL+YyHuNdV9D
L99HO7gR++06UV3QeyAyJO/DYtUc/gjkiB4mY/VtpLPicMCFsygnC/esbIuZIvJtNIgiSRkkEpyO
xgooH3hW0QYxZtEIUEIJY51MqiXivO1mjCYdCvWTIjMHCbm3aC9ejIt7tX/lqZP99YTLzEmljHFZ
R/RgNRDYK9X4V7nWTbi630BoMhbgXbJ2NDF9CnpTqtXFQsnCemjqJ9vkrW25VhAE/rE8Fd4F1pbO
hxWG5kVKVVV1PB6JX/eoMP1XLdws6Bbou6DxPlONdjpNbI/9i6tp1Iv5/T/UJW6yZ31pUxNGIRx7
tMQmRssqjJLIuncWsMD22gXonUoDZ4WQLQtac6sRiKsH6P4YQH56O6fztcSLLRvRoZlGHaEwUAZ7
GFN7rnkmFWxsKNDRltlRra1Jz8u3B5nnNggQVlxKna28yxRI/69AJznB8EdgURfSI+a+1wuhAdEe
Im0QuUoiBY5UXhutWxiWCeXB1qU6iUupTxEGTLt3T78xcLkNZFhnsKwsJ3AEmJ0idYnKOLz8xLa4
3CJ1b21UgfLhl9BZK7xEcrtMCTXkVut4xBPGCLlVVjdqvYk8sTxXyRd8Ns/C3GpwQoV+l660zZ2G
9EXl6BX6t01d76i7/sEEkfa3ZxCR7QC96YEMuR7jXIByB1cxrPZYESS7Lj5uxyyi8RzN7C1ZvZRj
O56PuKptGWZe9dc3/nfmp8sMxhoMhgx97F9h7afvpDhdDO04v5SbnB2uA8OCMpLSg3CruqBt+N39
qax1nyrAkbwLV7A/vAtIus9s7Muyn1smVF8RQJ5Qqa08LOOMWxmprea0r34Y8WN5/255fgdO7xLy
P9vBwNzRyR3dIpDOsZBj2qfGcn0NSwpcVrfonxtTQK+8hox5mqX/dL+AJyOG9VWNX1ludCMjFnoX
IM0knHRJnsrjZ2xO760yVkr+7S4BtDV/MpNLJvVGd6nwxlZcBd1trpf+gf9xfIIuTF9oeBrqK+J1
sqb1KqhcjNUow9F1PJVJT9sq0K9Go55d4UXuKrd1apQHE2TKgrQ5uV2DlS26KKwlMk66TEz50b4z
1YbVnRgoU6lANqj2orS1BJABGmqCoG+au+Tb5yNT+r6q3ztfv5pz+KoETLKW6xKX2mdq+UrfCyG1
l+uaVk+mYWe6X5pCL4LOkHS5ZeHGD12j63hCIvcCcep2vV4D+Y/bHgu2EOQ1xFZSdQXjcxtk5VP9
E+/hqreOSXWbslabM3oqL9ZvmKJPS/WCXnIYhdvFUHVJ06lKH339yI+Ve4g3y2znQ1sugz3FwPD8
ffiLOmbruS5T/TpQLi3vpBvW5YOx5gq+L0NCeQzzbZMRmD33ELfsfkYru089obKXF1YJRYKa6kmj
Tsh7OO7vLPdipvscg1JBTL6qRU0uMhju/4wchPkXrI6hEcL5E6YMPYkaBHSAnQHpymEermemHm+d
9Qk7Xw9gQTci2nWsT5Aq/DlLptQc8IXYH1Ystl/RaioZAfGUETGFQb8rWA+BCg7iG4VxkoSHoHsC
WhreBk2k9hSpCFqWuVYkiLmC5R+b8oSkukF6jPfIkqAQLVbAkSz1EUdtSMhPEt2E2N6bcdUyerN2
WQVQz8PsnTTJVpo4G51ZDtj9n2xU6SS4Lz6VpElU+xcDaaDfVf+z15pH6SvJkhC9nPxhcsS33z7F
ALd9C+hWNENfBMLzYmI2r+IJqDwbDfzT92dxWMypkfWFtbrVIyE2RMu5MpI6b3hKQaqVz81/vMr0
2Lcr8Vp0CySBtI337I/vjpEfqBrNkXkGc6FXgQjgvsxLw4VTTEzPpeLK/XwVx1hz8RUj9j/yhdDr
kUy5x8mUbt+BDLF5h31FocBcRipyz6mWSTjBzk4TjP1A1t++ZOtL3Mfgcz2cHRrujYuC6ryym4ec
/ewqMeRgsiIhq5ZuaGYbeyqENXu0AeDeCZUfImZ/od4Npqcno3Wjf+Om4HymV1NcKMeaqm42rjai
SuTj2q3YTYGyPLNVxdWswgDUqPr9jPdHdDOmz2380juYiJsWSeP7xLhXIg3M/4Ihp3oyqdeLfhqF
QAlEEHTP5IcVBPZLPcr8biQ8DSCpC+YdSMZc9wVNt0cgxZvlc9L0sQ8E1bJj2SwiBu4JOJYHC6MQ
maa4PtoCWye8zbdVn1HGqpC864aPaJLmpCP4a496wj5yJawVY+82xUxXDhVDOQiK887HjELopPKs
Fs7P7BbpBglJk7mIMMzohbHWeCX9DnsMRviWnRziz+11WCn8r057WgTqJW1LwEhEsf4ECTKY/fON
WEO/1NPrjrEajSotMYC3AZ9w3v+RnFy08tO+/YKKy2hhXcCDIQW5a7car2IHvctcQkDAsPDTEULl
ws6d2O0oWums3uPB4sSAS0JBbnsIzIn8dXtoYPqZnuzuipeyqTLDHnEknU49iPIWdf1CFhPSdREG
j37rfY5iPKIuVhhk4HBaRFqfAWShYHNqSd7+6seslNf9AzRwUDSHq8uTxHWpSAupVQ2yQAwTnKnz
ukn+PuOdSfMn4gp24HfCOD5K0ZoAT5omY/KA0/VtHI8aPyicCVOxb38be6YCg0E3nWSxjHlzp1+T
St8fGCpCSX0AZ73ajf3LZRsZgM9UjIRqbemFRczAroa8MJOXbY9s9pTtO47n52gf3dwdA62RPSkZ
leSQO/jXjhP36xutuBs7Cxc5s2Hj36b9MlWk6BHwYTjj/2XVUw0RhiYgN6RJVbXFBSDYSwHy0cUb
SGKrntOnIju6oC3WyDrz4JJn1uE6e8jl6LYtTeWWTa1Ha32Lq6OMIVP5jFEGE0293iPqKvIMqiIM
SZz6Rp/sGXTjlPibkWfhVZQNNaUt3U+MycbEkdq2PUuhX0D0FccjrWzg02qN5CSjb8+nHxN80JI5
PLwuayqy/0yJoFBe0+fi817LxezXJvZr2019TD/JsE29do7wJm74O+YUXFkgEaeNs2FklX1lXvSi
sedsnB51qYooyyV/Wmp2uzE+EGV+lriSWuHYfVALac6P3AlID4/gdyf5M0QjUPBAQLLSTtPKOcHF
rECR0pklHSEvarTn63RvfL3h3o5pnonisNWQ7f936TUwgNtziQ6snHP7RJndPbZujGrkkrldlmjY
ZchbWV2cDy5ZPaywWO+4UuP+zryUTsSjBfIlXhFR4iVV62seG5ZZhuF6bEmkCvKjrUy8n0YJlg3z
iSldc8g3qsh0QDQTtS8NyqvTkY0lvzDkCZjUbD+NBxNWiuuuIfnR9BzEJcRSCZN++VmrJwT2Mq6J
mftlEAk+xt2xE/ksX/AvklXxPin7OLJQefmdDjUx9+qZSWCKUWKj+GWsB8KoY1CS7dVax9g56/Qk
amfEPB+W7iMJWBjKMU8kXiAuaVKzSqv8D0bQch53CC50RJDf08ocJ9MDIUZ9I9V7ly7ob+QtlPzv
zvphORs2DHtL56uKGo9pqx2tyq3mpk+zZCZs2XxTGa/zDet5FC6a7jp7gKul+xPdPfIFa1RsF6br
sf5yl9zVY/XlMHXXejhZq0CMNJeIoGMG5DKc1JHC9wnkCQNHf0sPkx95ehvvzENG7HdXn63Nw2Gb
zpE9/98ZLBETznSx4w6nNFeI6HWwBcOlaA8Lw+IczQ2G1lsOXzZ4wU8D0qCb1ajNeOVQ17vUIC0S
yNoV/cjXwIRk1ZpQ+zCMSnY0EuVksszvqhJPEO7Qe/+mK7evdzITDKAjLmMvxReGwIGSb9eNzNIA
ar2GWFcOzKRTE1egQtUhOGKETnr9+WXU9VJbX/CfMc821EsH0SmWTjfp4VLf5Uz9dfct7jebu/1E
+Ve0/7teQ6nzzgJin211JWtsUhKfVVCU1t9yxwX3413ZMJFvOON+bXCBdxYoKLC7K96PY3SjXUFr
rjBQwp78yqUNPAXNIfTxjPKEr5v9CsZgOTKiZdAu/a4RNrP0E/iFTYAhlhafNKlzMI3ZgFab3lxW
umeK3reY53aGB8bAIhYZo3hpxO2VPtbNFM5eUeYEUhKHa55WvtK8FuuOdlu/kAUhHYKVTPac7j2K
Kz8aQlhWLuNE0NLUOGApuDZBwDFNU8Sa1IspaIF0mjyIlAKIDoiiQrOH3RpYLcsgboj6gQjuEnnQ
yJWq6TC54N4sZBknapX4kTuHQIYCRmgpb2mkoDZifeu1Oa0K5SuX+0jqzjEHF8b/nRN1AePOPBrL
UBNHaUYvhHNhgZY286imo+cv/nxjKOMS+5mXnRkqdrBhuSmdfZjLryZN32NzFQc3GTqEkrg5/gV8
ZQB2d0+oRJ8iOiB20ZFt+2MCcKgkAoEA7gR08Q/w1hd2wpvjrdZaBZqsvhkf8IoCwWKxSvKkZubg
bFQI3o6gXFXpj9PAS6c6MmRQSjRGsoLXf2yvDZBAOeNK3GGV2Zs4wvM4weGLmWaWI2x75jseQqDu
dlc0BUi4UZJTSxgb/Ful0soEyAjQ88G8Y2Zh0dzhu/3KS1xTumFmEgYr
`protect end_protected
