`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W/OUm8nxO3MQ19LHcqGZzPLRMKqH4GBnFUO/k8LYNBUY1hHdmQgmUUeQ12mO5b0i+keXJulmUxRT
qDEVuzXp4g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AX/Hu1HjEpY8YTkS9U8V2Yl9z9avW0fcLbUhRyMLm96vAxJsy8PF14TptcHRpDQ8EA6C14KE7UkN
pDGc2AHurZSiWAndag00BVuLzUah3PXkdSOnIKOD2rbYk3LumIuk/9SA+VCmxqMSHB8kNM8yms8G
/8YdkW4YYXoJ6wKlZpE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MMQOqWVSwcVzJzS0jIYlykOA5qcBdkP3o5smF4mNkbvjhXfNrbNhY6kaos6dDPr9mu8+xtwQFCDP
gWy7V86AenJ00mhkgIYZzblRTu/PkIL1CFMmyA7xuWPASaF7SshvQADa4Dzn+MqVKp6DosLyVCaj
+pjB6CnvN99G/nZaPzAmiqjbN3gYHD+DX4Fw0xzWUYW3gOV2+WQCpoW2tB3XRVk3U/hL44zOd76C
mYyw/GG+Z4dKTOm1n5EiTaAyOXdeRUSCK5KEDiqZCJbeP3KcLQNPxCo1iOuV32jjZrkbS+IfhniC
afk9xpTD8CbcqZ3XvY7jDCfUHzBh8vfiACDgQQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4Zzi3OqlcDaSO/45uobjo/c0tklK/qtoMsDK4JWp+EiNICjXn2hJFNbVnNoDqbNOlbFZwccMwmI/
qSoDYg8WyV+Ia5P/ZADnIqu5T1JhkppW3209DCxMr+Qmxj1BZCqS3xp2Zo46ALsbrQQ5IT9eqHzQ
ozCyROPlEa0MHz3S16Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dR/Y0crU61aC5qCEQzojPbFvADNVZpBmMj85SLiBXLDOnzDNKexNjcecLWRmMJrjsHn5q7TQNE7B
GicaNCFAe3I+UBm9oNEPJw6qDb51B+oSWv+JTKslRVElrxKKahHVy+YWHe6ggtsrJ3hZfTxs2dpP
2K4J98u8XJI5vaVDisPptgLs66kpP3CZQSuMB7mvWtobl+oLmTuV4L0QP8ptMF2QaSBEuKhJThyd
fLZJcHBX+U4DlCElS3tWAr6wn5O91IyuiNNbRk7Efn+Y6J6pu/Yq4CM+hTeSgi5jfCRyW106wqJ9
ZMT+GGq2BwyPpbgUSRlljzLoZ1KUcZXKMwA6Eg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q1FB7SE26Z409w2uY52ldW2/oOB6flFPNDEHcy/HrfqmkUwovMyNAidaNe6+TosZtcDGRIewIJgr
hFDJy+EUxK1VjSJXtvewu0vZ87J/dttgKOCRkVNTEkdIjgJzk/2H2bxfCMQAHcOWIBWI3RQ7sXSM
OcCez62kn50rsNU/CPmHFml1hwbjDGqPH9qFNxEjxfqmJezJbkMRq1qJIXSasniFUE4U877Uigi7
EnaBeWq3q0xemSwS3sSuZtFcGPInkBFt+STMTyEjzlo4EuAm6bUcHDh2oHbJGSb/e12U4x1r/t8H
A/cYOghbCnxKPVFV3WoNCmNSU5x29fZS52sc+w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5392)
`protect data_block
ULDd0RQ2E4HpVxAXpJYXiMijQ/gny6Af4Qk2uyipVjY6gT7FbjMkLKPYzmqdUXvy5dsdmel8QraE
PHJOJGLxk/2pW6x3KYhyWSuJNVZcxMD7icITLadCOjhwQ0OVs06sb/FkFuz5LTKVlFtHXgB/WLGT
hV8/s5Itumfbtr81A3h+VGxcJHOZxWd/h+EEAhNMwvI97AF7wLf1c/oShzTH9IM7XqGxRK50REOY
rcElFOphMjWiza51PIm5ITzP4yoWFJ20tqs9OFqwPgd2uxrIsMtbzSFi00AKluAr6C8tNViS6Q01
v7LnoOJ0xxz7JmE8RkiqUs87PeacItEhiQgu8c7/snL+A+KeEsfGJymkiyYD2zFuJXKkCflLJA9z
3u38EuzO/TnfMvlEdWZDm5meo7qFvTLhwoB+WdDH7KhvwvTSNv5W7mvgv/a/3MbeHkXSgX0QMXjP
9qyZr+4HjxsnRK0PDBIudEzCRLVgqcE5AB/mcPxRG0bsj2lpZsY/jBc9CIAdP8vIM7idJRh6Zolz
mgLAti5kdgYM5mki/oQIhcc7o3DfsZLNKzFq12JQG80Wf0UB3+RtM2iuvgjR36OHy3fgfa/yvfnF
4rH9gluJDPJAAFqSvnhT6BDCWjK1raAtCHRLPDAGNenxHbX2W9L28a70gH2OXMRmUmYm+Z0xL8p2
WVxSL2ExyaHTN7ZL2yTroZO9Q49r/kajMjpkyQirARZZsLIG05ZVygYLPko3o+k8xEjnPNGYw16K
z4yrlHj8X9oXQWN0skQrvcfDQFKw6TAEq1tPpINrPYmuvnyhBLh8cZZyWXEUgE3fgtUjtnlFvA52
aceM+MHGkhZ9uoQTIPV8Duyh+QviSxT9u39xVDnlw8VYyGwWxYnrPbx7/6uG53RSzTC1ewT7w+BW
/BFAvIbQOyPLGdjHeYgMcWK7ZaemugpYZkyJlmiIfob4r5ZqFfFjvtp5+Jra/FlgquM21t1Dl3s5
wJ263ER9W29Fqlu7Vsd6mkCkT07+cgYT3/dv5FkfhtPH5IsOPkFfAsRnoTYtVqkG7HwaAKGNePvh
DRDdHPLs0kq7LCXQxLtSm3JiIdT0ICItoe8B0RU4VGje7FI7Q/+pLMxng7xwBj+x4Zrps5ZoGplL
TOH4AYBlRWdXi3z+kdnwrfqCQxhJkYp2ZwtmGIwNrg0QC2YJdC9U9lbnbXXoOxiDf5i3TJpaV3uq
kqY4SNLf2iMspU12/SDfx5fGm3vkkf0ko6/fssDmIBLljBLKFdIlihwjC9dCr9WxczCCFjThLZtB
+rvTgHlA/Ki+5I4cy4Jn0vPB1MxXJ74gFEq5qFAyidXxTJyTSG1AzshDEST4d/bN1hhQnIy4+iqN
4lRbSIjJqYM7851YBzGwPkqQ0Magda48tcGd35JtRbg7kKOiYyWEaiJ/rhV12cnIxi2JNlXnBCaL
5yUkbis1VKm2+LIiFKNqaRb3kV3O1CswO/EpPyv8pc5y+BGZe64IFRDaPY0XZAXqlgHcxcZ4sDZX
lYSvaNsBbcBybn4nTqIVFYiQnXG3F0NobOOI3kzNGcHwnLxOsDQUnEGQpRy8pJG77E34cofE7Wva
Luulnr+tOLIIsgWDsea/dBYX8drVE7T6o0mHRrbwTP4UILBdvGTOysS/yfSYE0+PvcrHbqWfI+43
oyuKlxa+GQHdTkxuQqdEX32/yD/Vc0HgLNW0LOWGddZHj/yGc5D4oTf6xph/2kOvaOlwHMSM9Axe
1BQNeK+pTTmJO9ySE9ZMID3KUUi+MZr4BpS++rKj+M1OiiBJg8EUGU/VwZhPSCx3JZL5GX1C2FOs
LcqqmFltndi1eaEwVY06hBMetarejkjoq55pyurWvu7PhgATclsAgcDYkatzmfIi3mElE7dOwJXH
qwFx03C/g1EHrKsTrXDL0b2z5FMbZKTk1lAuhYQrKH9ZcgKNdulccfdONu01F7ACdzJevtQ1wE6P
jOEc6ctOsMGD24jbWCjcxbm8sy7Tzbv5MddU6I61Ti1avFI60Rrhr2fDghDE/cI6saw7i+8A7QVX
7Xb13jBUYfil1bJGQ1nPuCfz/lM6SbngeYnaRKw+tj1rKIJzfWtiywwsLH57xdR+eM+iIxTnz/XH
jYEzfstLCuqVvnLBE6TUYdz9jD6/7+7OLJRLuewjjCOUwWCakvPPlWP/J0Rt2cH9FMvTLQ6/IIIP
diq3YjGxZRRoZH2ZwEiprddyiAYhHOPembIk3ADV7pmfBzZ3LHqbD9OcPqAXTNnbh7PFjIuFWMQy
r1pybe09twdhBNbASYKHEQCqUX0bhczAjhWMsLsJuItGC5eUQFNLXe1zz0ZhtkTLa2249IPfPXXZ
TiZhBaJM7V4zYYg99J0xUnVvAd5h/J3Pqx1/TgmGSk6kT9Z58iAWkVxe1+K9su2Jch3lNxkHx8PN
AxOhk6+bm4vn2LzxoSzCbaOGTBtSRXsVZGuQrDEsj5AHscDGCqeVczq8+y/Wy9YOHrJlSlQ5QBQK
iCrRMfQRGWIEiVmuqDm4vQikkPvkRNxZlEwWwwhJa1JCpNrHpQDrOOg32Lk7YXl4kP7TdB4ivowP
bbgXSIcL3+vKeCTOGJNoCrbPq1YY2senMyVtk8Eyva1jq5uyL5t0A6KaukWoP0bDFmk5wuCvhSxw
tSdxHk65iHCUhfb8SSxSczS3xAb1BQMA06HQCMTHWG6maP7hs2Fy7zeqSkCnRQpdeHmOCTa+06+e
wnwjBnrB5Qkck4WL+LDXk7iosY4MCgJB9I6SQnBu8ueOkUHgDKgZXJudEFhZ0S4t9WgHl/5dHLRw
MHBHJx09hQbZaJlgc+otJevd2E853axcxe3L4xnwljE0jI02HhZBGwuOZGroGc0Lp/tve2Dx45eG
427ne6FLnkugtay60T9Los6Mr0fX0aJBVPEXS1FOPj2T5muGTH30OuZfFBUklGt+tvXASP/+byjs
bpMIPaHXCG46i/ovIjZVM7uFU2stn2pNJAtG/5oETL3nh6J9HBdvCsFhaTdq7pYa3YNi8lJi/uhB
P2ERzsojnT4eHUPVOVgvOId3kg9zM6lo36dg60kKePTi6tUc5a2QsGF42hm9t5cOUeUdYaNtLGTM
4zjBrGQDykdHxXTi56cjRgg1/nu64kQrSLd0UbVTQSkr8EQUciSG6ycPpPhVvqp9Fn05sUwypZCS
cHfBkdACFI6X/Y8wU2RJylmyVQXitvtOSusymmaagoMSJLgk7Pb+IRnuKsVtPBRCcU+ReDLZf6dF
fw7A5BdzWMqg/7SHbz+TNeoxzWpCMYznYebQhmdo66iweH77Y1YP1WilAcoK+z4Idrri6uLXeMyq
UiDZOBNzD064PS5+Q2pUYqQeKP4jM8X0qT5LaI5lpAoWsZ9Ra4QHw31n0VyI4nzTfGyc6G+ZDnML
mt48UGHisuCkJxkCznepuhoZGA3FrQiyWh+A/t77W6crG9lmIVRxVq9txs5Ju7sO8oASB4dm9+OA
G5jq9UUICbmatc2iNSC+NEQfvNyz1WxYsBL7cPf2Wdc6XGkv1rsFIx3JTfEeAbfo01INwSeMwdyL
uT3dle+j2dWpSIl+3CpfLJHPSfdfT6GQaILhTQBxw/LLVxGbX7sSr4mGjp1ywzdv1vq1jFfF6Or3
cYtgn/1jtiNf2Xsc5yYMs5LLDxyt5trsZK5CWOO3SivwVUSlCtajYW/GS1T/2gtJKEYMPMY5g1KL
k3uAm5TmedQAU6VUdFi9FMkvoLXu9ar+xNvEtj1F+GdTk3QZO41XiNgJQRblH30kCeJpGRNhoc9H
AhexDOVQdxJEwe9FsFRBzl2m4/ouOzPgoGVfO/jOEKVrj84yUfDDgLNYRBLSr+/UIyRZR5Ms5zU6
dGQemvJfwWoNiBD4+1QTfspQuDj2pEXISOTJSuUqtou3roZk1QiQ930hGtz4/f0Vwh1cgjlp3CFk
YpgmvK/q8z/ylxFrlsI5AFJlzt2Pb8ybkR1RkKDRbBPxl4KnO8X2HCXQssSlUnkG2hZcrxtMkqKF
/Fl15k/bNXeoDoPVbeJBdJZNV0z4BJTyy9ulQWBxivWZesn22pFaRTRRTRE2sSOGNSeCahcA3v/+
f2k1LG3+JwjB27RLK3YX2cbXlgXuq1Yk4I+gO4xUTn+Mph5Y6J1YYmDJ0Qn53EeZKmh9g5IgCnV6
RliU9h/5nAcqETXxfLcqh150jize4dzIbo5UloDQkqFLTW07CWSj4lAev5RQPmRnvNzE6iYvxz1Z
wpbD8XynPbtD9r7OA5Y3uJrNs6HPiDJIHFKlSuojKiohW0pAAFwu3uKBlscpA5TwoxWDURmNjU9o
49T/df+6gQ1aK85dZdsvMDGioa4WPkbRscqfKzIfykgT2o9NAz7IUW+4zo1G7NRx3skl4Hr2XwOz
e4bMLzdJxWXyPIesPqLhPqVlifLHUK+/jTzDPOD7SGFLIR9MiKIYp7usvfgOvzUkMFNuxo9cdufk
YfuCnCn3LoJyV6Ha1L4nhR14Ws0JD0T6PmqMSWOyjcqxo3gY643sWVwsR4f4+uiw4duvfL8MIEf+
4cJK6/mbUe3s1j5UKFfA9NYamj06xPjX6JTIVLMsY6m6neggi6vh/Os++BYlyNbnkWhStQM3Iuro
CWRZlUF2tQG3jVlmZJY8HuEMlCO8aRA2QdU+PXNolyf2XFDYoLkMfUZRmzj+Y/tucYQVTmYusTkp
x67hLeuM1cLZxz95ZR9nBBUV3r1sQGDm95dNPylHqfBBB/XZuogmgCewqX8QAi4qs3uGzNQZWSHK
mBjVXyKqW4LUSgMbvNd+qfCYbOOvXPkuziIxBE+H17jcKQPcVHrhiGOTXSdARoZ3NgHpAswjIcFO
1/iejrdsiNWHHGk5PO62kB1IUDIJddUxocKer6pdX11N4Qj5RRhE60d2xSI2PO9cPHeUFYJIJQw8
Zwcr/VCicgmF8czVg3XKCC64fq+tD/PhMa0yaYd0GHUEaAYfJ47zDqY0tN7gQuvi8dxUHMjBsPcd
xm1WdY8793ZfZCtToWJecwRkyfW4Ydyg0tEou5V55nv0xUPD5jEsHbCNKJcveRbAZ918B77bA6Su
dxJ8HuYYn1zrtgINR0PeJdQ+W5Gi76MuaiHKdPOMh2LkYAg4BRRRXkzPAWLbyAxH8YFzFWgYjP1B
QaXAYqH6DwZv9RkUWZnSFm8x54P8lthLgft4NFJEZfA8e3I6FroSHj+XTcp8KR4NnGTkWHKF1dwv
Lnv5liUtK2CT0xakfarMxYgepDC1ls0Y2GXls43YsRkCDFbVlG6SeeEy79BVTit2gzOXlMmnCmGI
jWuu7QhOqXxtY8WzJaq3eld4RS+ag2gz0K1vWv7sAXihHcZv0f0vCWvdxnrQzlgFjY3F+k7Sk+YB
U02WGdz4es7BVV66Zlh8vi/mq/cee5bkfHZ1gLWoH53fAgSWQmmokzZm0wExIgmAfcdYj1c5NP+q
Q6fOV9XSho3hcm8AtINQc8UekNhgi9WMMQeAbLp//gFpqB1kKuqG+SQGZMrYC2713vkmg5S0xsRC
vT6dSf4kVTqRCPc1ks6JcnRm2iMHypWqxB0aWWgYb3F/bCbi0gM6fU4n2ignxpFyJrlegEU/g8Uh
fzkfuu2FMBWp4qa+lQxoEjVEBu72wYrk40TG1v5vAIswmUnXGlpUgQrtAaLaRZK5NtKdDyrHvr0k
1O7zf+HDjQcDDTZdJEtt/47cEzhzXk/Ctf/0ZfSiWXQXIBHuk/u1ke3ex2YeeRM8Bekt7YArQYDC
0HdvjeeblP4Om4gR1pumpVSqPjtSdZbV4wXWaFfqo5pBqlxBDx/VW9VdmlDY8X1Db/xHHxn0owio
ch1PBr4V3hD3IWIH59ySrQb2wZjYR7Mqc4lpcGII6HvW9dBHWP8T2Is8/FKJ5zT+qAT1Yxlh+n3u
XsqtlJgXpNLjDXeAUVXg82Tlh4aq8tKmMVMmf7qtULuIoCr0GtUQ0r1oBWCc7Wl1bTJrronbHlAX
YfQeDb313+K0bjpDp7+9LEl7/3X60GdB7ILebqxZBvOZ6heL6QwMDZGroHKCQ7vCI3kG1m5ue3ZL
esPFVkQYTUETd+99TAZ7Q5+JvCkl7QG3h8V7uGU4POOxyVwUoDqCxijnWVT+ee5w4jXyBB7mMFbb
Kp0rMRaiTLSmhtcypXG15bPc5f9L9ksP3QLotRFi5knuWbF9TfK0MONR1NldmHrx3nzhxVmHIlhk
MKrlEsLGhFO+FVSoXaVMEpMBoW5eMoGRn7ggUKc1D9icjAikNz1PnN75iLXLtyHiWz+k/f2B2EZL
dY9yNRqHP0nCYVSlRdsCb6/S6Ne7fOLW/GOyardz5MEE07U5+idRfGcWxksHZuji1CsdeSZA+Qyw
LTqfdcUmLhKKuOfiX+VIls/QJFCGUO/lSfuwlBMx9QJK7KxPjrtgMeVSFnPEkzf3qKDskA8KROLf
pi41hR2Q0+qjGq6BfTvb6OSQK4OWk/QcADyj0PGDtoiOKZZMnd4drVZR4V6mNbuBB8rw5EmmoWUA
W6MCLl0nUhRnPmwoPu6Is5v1oDG/dDqIVfh0jBqpg4YNCe52osA5QiLwmnfwq0kRZQqRCMcWHwn5
v1I6IfvelCCmYeIMorM4iMUmPgxlBQR0JutYgCuhCFMxz4pH34hfWlmDdNCHcVBx/wYabf/3uqYS
zPD5c6pj1Amy1A74vjNnbBSXawbwYLWs01pRV9fsbrgaO9tncT+sv3IFcaupH0ssIRTCMF3tqUBM
r56Lad1rp+B/5ZAAPfw1VIx75bS4QJHbizvHfFSZu7NE+n3nU0sRtIr7Iv8G4Miwhju3CgYyVc8Q
LW/NYUPfvZS3eXsgCQALIsLh4Ln2vk6TPOKAQtJkU1nVDeGGihScEE07oH+Zow6vtA+APL1WpFVz
CLmm2q9knR2997EK9bPsU3GOMvDZslLAtGzav+9ovdM0W7TR6ldTj+1di7p9HCm7cPoBgIh2Q6hq
kTmdl7fffrvlGZRneSTo2hQHBzKTqEGm+0fEY6+fhe9YnS6vy18zoXhkIVFsbRHo9bVjofLkLqv/
j1RY+Y2zDP0+m7vYlei4FNvrlfP3SbcoCc9KKNLFK+Vy1o3reIePkc7+A2JrvBu3hUH2Nz1oqTs4
ole8suV0HznLaLvsKjvmr1Tn9UL1/apd6Le5JHzV7KgUMg==
`protect end_protected
