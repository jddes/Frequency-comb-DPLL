`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HXsCLlO+mhER6999UqPguhOSLyphOCAPWGYV5jW/TUlcrzl79bHLUR4wDSf2HMuTSPCMzf1gBipT
NCNdtj0VVQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
femSaA6afEiUsIo+AmOu1hAlf9T4wjI3xmVCwthfqlHWHDkN2MjX6Y+WB3Lb9nowNnDsdtkI0BiW
li/6nDJWBGQCbSYXX2lDLotUz8Fx0tltxXJxdiaWtVRK9Ww0oOXe4fDwFjmlW3CLRb3Cn/+oVsLT
tfypXTVMPCfoHv6/uMk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ssjpHcUCaAe6fiO/ZAsTolYXiZ/vZYZL5+dG++I0tC6thImrQ8Afacd/RV0RWzDlxYhGAOlYFIqZ
ccb2jr0vJ8k222QtzNA2HagpDsqVDO8G6DEOV34nk5Q9GRw0fphVrXlLYgkdcB5MPZ2z3hbbztPV
khp6FkenHqXf5xYl9jICU/dWu8slpuqpvUEt6640tUV0wU5/9o0lGTTxtRL3MMb91w+yq/AniGTi
UXHQ1PvVIDWKi4qWUlCh2oxe/46XTwyk3KG/TiZcxNxKiKctVme2prqAeKinRGi8hTBke7ivNU0z
SBgjTPo907ZxyR9gbWrYSWSW8wdpDXEzjXz+Hw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CJnz28couMgExB7wcn21QRUd41AMjm0GWR9Qm3JugHnwVYBIOFiAy4Hulw6I/J5XNmcueLBdEyFu
ug6xgEXaLTTJ3r8VGS2FQQOdZ0ejdbtUAiNU/NTYcnOSIdWvowPsHC2Eq9bbfNRDxW1KqIgJTmYh
V6GmOR+5hL+ytCLh0FU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p/oh2dN+109zc0PJ5NUnowr4V2TRN7XOK0VeaCnPeewv47iW/31lyy+Y0mBgYaDlZHfzDFSVWhf6
AIJbuUuBBSbKWY9w/Mq3gC95OJn5Od5keesiv+RDbOeUwisST0BQZGVgfn7sa3boPGTF5mTVn+/A
sFrYn4Ue73mFTl2joA2zGSAS9C3NMF3MzB8LuTAW3VI/2bc9bR7r9f9ri13lHAZ+Bo8Pdymnqcnm
x/2TdaUZudgoFmXOOArzUfS5IzjmhZT7JJz1OVxiBhBaMqdQ02lVlPldOmE3o9XUcBfHASzhACdV
IUhZA/7SFxJ6S5u2WzURAyOui49JQ0/CnwLLiw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
txP3I/W8eJa8dVzaHd+kQNTcDDXBSc+QdWRpp84GORUdckWeIJPFU/fN2i6LfaB7NzVdnhqaeDB9
KTpgoBL6R3fMOwiZwsqtqtpRE7te8IqjbgHOc7J0pSZSEhXuXjAnmfuZnwXw2Bo32ZmqAsJkwwnI
lnGvgs86jo2DdoxOCLLOC7Mgz0povdeZ3JZLeP7LYrbgIOSQV2HtO3NFwtmZaZCFlXUzf+5+UTzX
CqtjBAh09HxKU5ICzZwBABoFatzi7BuvMJFhppCKRWtgkvoE/1skYVklMW3PriyjHFSCxTstO/3J
mr64n5jMZM/1mK8jaj7m7X1u31jLr947qxbdbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18016)
`protect data_block
G0h0v6QdkwBrAAAAAAAAAHakHwPytFGCaCd0qrT7g3KlH+dw0xKrLW+C6nQyjfDDa0Flh8kF22bP
AHKQZ/8XnpK4yClMgCkcQF6J0Iq0gOX4TZQG8GHpswuYjNlO/IODi3HqpSft4UKaB2Pp7+vK1XNG
o0dqblIc2daXyNRZ1iIIeU29meWhf99YRIVPCdbOgnr7bRm4SXiskbEVkejBaFLIGgMV1dk0g8I/
ZYTpZN1kH4yK/lbVTBY6xQzQ2HweqMFCnigVhnOa89s7aFf41NMMtLb0oicVT6G/Zk0JOrCLJLi1
dv7LrIE3EKTCzyKWvhA40yXndmGOXr2xUZtIwWEsKGR/7+rUSXqpdKixAD+I+ksnmXVznJiNbjLJ
hV9hT3iMjvqfOnVUhRJG8JboxvHyXsIBE2Ul3SSMtKrdAFbD8UapyY8r53M1AO+N6EFAy7WiD4dR
tOW7nLeng6oejv8oyLobQ9JUZSmmENcSBqx7aW8V+SPEzLy3Y++44vd65aHgOtOgqiR59aSvnDOF
qFpnbGmuQ5hiajGCeYePF5lqFS4C+AOLzt21jw7YUn6K2zElWIxzBtPlFngH94bauKZAkInuCo0y
jNj1R+/E7Tud991dMOmaKAGwmUC8t0nDdHb2LX/bd5Nj65wlddKzof6vZ/ujzGiazhiZT+kq7d0e
UWhGECCW5KJWmfxL5dBCiCsYbUvaNQesz54M60IntHMjWbhMFsukZwrUVlgigIJ7MqoHYcU4AH2b
T+dAorSR1pQUyqvMmaKosf/jtq55khFioJOHfiVng7SxscnhUWwDrE8CW5hlyGipHZOiYxwtf0NZ
5J7s1iDEJzpLlLMC4m7L3Hc6RSAGUlbfTRayckcazi6Kj6DDv34Eskl6bx/zqAItQr6BLwcuoT2d
8NSi07jo3fii+ca6V2k2GK6HnltPbcnteB2Ubi6FH9uKRlPw45r61kY+mytfr/MmD8C012E1IUIp
7t/oMJxkR1G+tL3pRU8VXGc8aquZ7E2X3LDasxukW/ao0y3FROzsGlEQQVAxt98B+2/dhR+c3GPc
br64johU8FIV5rlfomO5tMX6ImID/E9nIy5Wv5zW90W6Y4Q7bXB6U1y7KP5sEwkpm8WVl3QJxVve
EC4X3POa+PD6uy61NW66ZyEhOjO0b5JAYoAg6MJ34GawfM6c/e0yny3lOfP8weSAUUY+OJiTCIKb
PujWZZsnZhjUddBzNItcMpvswsAHicAFzNdnhtX2C4GfWFuEiLVrL2hzoEBZv8qv9KQIKQWn0s7o
fkbJAIx5Eds+KzHlwmoFMZny+rLK2HdY62VNErwuZmYD8Ov8p7Kdv0K9TZt0tPvJh4mGkAV3edA/
56EdaJOyby3GIaPTpGxrqoujCzimeJ+ELf47EhgkCRIr5+CHmwjwdxOAKUz2kcdj9K8DPuZ4zcNO
hO/enX+zOj+NicA3FuXk96AXtcIzyeRK6roIDkUjAkw+GM5S2XadX+98RR2QX5wBDgBQjkWYVfIU
PMn7jkgEMY2ykdT8hNYi7ZF7ELdmi+5zOrHarzRAuj/T2IQe3fmOB0JWyq6iFidt2plMpCSZszPh
nI62Q7WO7D4Yn4KqoOb3RfZ3Z2m28OB9GDNGttU6a9qsMbaSuu+gIXWCdBjB7FIqAtaRYWX7MiMa
WcIFlHE5L77UYisk+E3C8Uq9aUUmpQzIUVA292N4W+t85JNBts21GwCvhe/Jima9vKvgd0nqNCVV
sIcLh/CG1YImd0tMnqxiOuGFmySLwD/mAQWL+BExI9+dKXjNhEZlZNW68xdOog6OQqXTWHWcoANX
mJxsrfrMfOb/d8xda27CrBqkLB4ipJSY/kGKgF8tNRd+gyYNoMiaysF4j4cZOuwJLW4yzkEo+Idf
nGz3RyMDlpi/q/NkQkj+gsQ08PTicxiF9lhbjDJxcaXnuCaWOoChVFg5VLJs12xiTFt9kMb9hcpX
GqbrmBjyOFzDQ1A+LmjASZbfyOqsuHYULUhkSd8SbuT+HKamOH4LDUPWMg7XTS7dOmjS/fdlokfL
Sp98upzCNWQkWIicBJdg5zRjEvLZuR2C5kh5w0ZbHFCz2+MRq/FLdQJc1dAIBwx8bAB8u4Xt0cu3
tEYLXPdRdyoZOA52ftT11TWcvRH/fN2UZ7YkkeVBaOtrWsGqB6yfUKOd0e48438TSK52aid4OxvS
9C+433GMk2++YvlPSPvje1tCX2m81QgAHkouZvmGeSYMDFd8+pzSNGOeLmJfE9eZj5Y4mRU7vHF0
xCVNp4vIQwj/fdMz5au6aVyYLQPCtKkIl+PnUI4wt8npMVZ0gOCMkd35wTSREhYtWXtdwUdrdYZc
VTqpYkHunILeMCaJUnbZubl1d617O5hy13jHeUGpEj+vh1Dcje8hftoSdkd8IeltBdN9/6pyFqrC
GpCnHUAhtFZ1zlhaFSkqevhbhcDU7SENpViSMi7K2D0YHqVimo2w+XgSah1Op+B1BGhyfpE+/Xdj
3VthLloKWIhdFnl9A6VpI82J7gxModFPh+riNc3ZYUcXQ5mLk8ZUheQnsgWKRwA9vSo0+AqSRSfQ
Sr+v6+UfpZlgFnCVqZxMjAz27PK3PjnAJtW7eqE4L5v2tBnhnR8KnmRBP+n+0UX0Jthfto5m8X5v
9Hy4z9r4PjEwB1um2E9nK7ezd11iW6wdUT/b2N/SkwecRlejKRvzNJowc9t1Bp8WuubdMyxELcsQ
CsG9lK03WoOmXUEVlmq0bfeMvf7i9uc7Y+2VnCbhSAxXGPejJFJOi68Qqyebv98AQ9iAzS4LOPxW
keSHNhn6yZdvOIPCWyKvnI+xBcxSOGTiiH13F7ZdOrIWGaVkQsL3mSLIdNfB34AJW0yha9dpfrTb
T0yLmgFdYPlHeSPsqJu3vi+vi7UGCcjRMtPSp9hcpjM+zyFSTyiHcmZaEGEex8Cx3Of8Gq5hUgWd
58ZEzYcYUG+cGGRGi72jqzKCMkwCnhFFcE1A00bzUXwlTkTN919KLMqtZCQWYVjjoJGuNU+d5Mxd
dXE5wNJrmYYz+IjVq7pyTkyyXUePW1AB9yUVhxgEmlQg7oj0xewB9eLVT9PONx3GTIyw5nGoCoBZ
Oc+rL4FtEUQdno+n5VOVwI5nQ8Gbx1f4hVDyvW88ZMPwy2jC20B1FCyRjEDj44vlCYNoHJ59iPJ8
0cZ4I9k7pKXU19cVBNF1oDxAGfqv1Yl8fcaEfpNXkH4o/JU5Hhjlz4vQoo6Pg4OAKNUKJzjdBXUl
9t+saeiKxKMvbXCbVtMFnmAJ6bzldEIFlVNQVe9eX0acxwQnhATxnYdoky3Rg/XeGv30cLrae2nz
jxRCJwXMXrF86GHAss87RzhtuQx8F+Zf6s68ijyvxXAmizB0ObNOh70JF3Z8h7WOseebcNoLv5xJ
puJ7groxXw6dHUqM5ObAuCcO2u8DfKoZPI6lNJPtUFFCCegzbulqduX4mafc8d+YrOSbF8pw7GJ4
hgGiGcYVKZc4XqgYeDa/jKUxtmLXQRKfGzaV1dPBnVppi9aV9ufogpwlQFPL/zDcCGaUQbIs+UPI
/UvWbGWoQoZyDr3d8O0KSjzF0bWj354iMgbF3IGysiopgfkMKACFAQ1poff8BQlWxzGaeg1hHIJM
cfFN6GS1Vctai+LQDsZRmO4mh/hwwR+GPcaYUdNcc5g43qpSKuQIn3ppSWk4lQxsgA+gLdEZz6kE
QrdLS4F60DtqgfLKRX7gjQ0axKXmCJSva+QXJVSaN0wiZdRpc04bGYVZnXh/NLkdBJWhmH9Ia7Ro
2sRwnH+iX0Avc0hK7wo7J1oObQylnLuz+fIk9no9UjKc0qRitCqDzklb8v44tdb7liDDRYCbW6jm
a/ULni9J6Km/7hDtYHGX4xWupcgnV38lvvlXv3ap7TaHbjnAWEEqtpgBDSxZH6tYCpworLhqhRjx
gMBj2unK+PFLVWw/UMS9X8K/UgIy3ZhkLmRY/AbLLF9QdoeFFpTN+m+/RTLD/srAQyLpX4U0YOEF
saUIvoc/SISTc3YUgKlwqSFCMawKNThfgJQfqBpn6ZW8G64izl/BVFz6yldyYAXBHVns/3ednWIL
CqYG1UVS6DR0m3in07edvzti/dbaWrHkSFbpy5bXN/WhiicOkUjDy9SU3g11IFP85TCocTEuuIcY
oorT5X4epczDytqwEqONdOTVpnY5f7pRQ19Qiw9QLoah/krroEX0AnVVa24dIFH9BZDzX8hYyyUY
NEfPe6M0VKmzd8/di7gP8/mxI+bSZr06DhWhjUzW72U6AUo+qkmFp0Q9+58dndJ+D9k9XkcwRho4
ZFVnDC8atElojFby78zQrhVZs+QsJm5uiJzvUvoydQGs1GN/fwoxSNVbuQ65TRxIsen26ZbmBQjm
F1Mhz5wx/p15gg6dXNPb+MscD6rGf8E5a4zY4yIBXZgl+//TQadtvbP6a0QVbuMmLxPTtFeuO7xc
uHHB4aQb6lzAJ+LKQGjztz/RxAyP/dkoEXXSA/ZhsNC4LBohupFxRFe1a1kyb+aJmJVSHXjRDxe4
gdz00lIHZejMD6FrHQ5iqFOfGA9EhQoxeF5zfXcQQoJwt1OV31ijzfMXfQLjLPrVxU2a+ptygTEj
ohVRW8cbrQkSpjrVfCjDpxjZc2JWi4EWQ4L7cMRq282TmVXI6y/wqU4IvNuGaiBj1WyGJn4ynaWJ
3GARUr6dqKUN1+utuJbSBrILpEVQwSM0FobX0uyDFrTigfX3TNma8I9Clbxfz6D3hYM3ec4XsEnW
+XaIGpiaJQHlJIvGwE17rQthYkqD16rJUhEf/q7VykUnafyksnX1iVNnIzeUJUf++TcTfBnBP/cQ
P+5+Nt4+FCPsSXem/PzrIMeVuS+RP/+FwcoVQBSpLOr86wPivojOZGYjRsAS0kRTYS/b5+qMNc7o
Z+RgNshp5kamuxw1NaEpVRkzNFWrXFqRPO2joueMqtAW9DQts4xIC+q7fpOEb+5abpVDnnAYf3jm
DKZR77OkCITHU8bqaX0WW4W1Lm/SExSvPtRQUS9sj519Bo7QEyNvK37v2joQHioC/6wuI/w8Ycn7
Zw46d5M5vO45PEUzqsOBqRBZQA/R6NNAH3zW6cCQH+oLHVtkK4Splrp4m5ysU+PkO7KRk9BK8JKW
8ctJ6k2PXFo2HaJfxNTjXtWpV2elg4JNXVCrXZ1gXOY+3kmy6UCXHaIvmw8+u2vrSXMG9SmqMll6
Gz2WcpS8PRnhfPuLkGm3cTYob7vbfp8QRNcTu+zvs5qRoPZugUJh2nH7Q9q4QDrdwv9RVHr+hQXs
LcRpKHruBdPHrUxmlKrKpc3lbJiEsnpGkO+FAuDU9LXL9Pu4SPCm7FZGlPb0GIINhWcS1QENWFWO
wKeMTOhRPe4p9E2ZD83eYDUt8aSnyhoJUfXADgXA8fEhYzvnlZ/ifEmuko3y9e471rnhxt8PsuEM
5TvggkbGSQFGI+DIUsCQWUJmc+6oke2H3PEO9D5Esu1/rVWtDy0jHNanLOhwb86WK6RwO6PNNZvy
md88X4YS8Tk8+lvaGPMInSVm8vl2j1GfH+JyDSmlZi/b4vQhOKKE269K/SjfB8y7pm5ZJVKEKBC/
2K3GtkwPKKyMWdMAkAyIWVJwcq1hZmxXexexn7ta5F7H3RL0YyMBbIZPL7DEo43jkCps1JByQIfc
KHmCYMjhiz+6H8zVLQA8skWJNNJkO9K2aBBDofHBTG2hWkL2nbrapCpH/fUnrgwPKRdfjLQfeFo7
ggbsk1wLYd/VvWi1dQZjjDL+ts+Sw0HBJPB+0WwzASh6iqyBaoFuXrR53kL8VWup2eJBOcNjpBvN
PPsm3/KDB9xlILcdFDpq7k5dlgJIPml2w7Bt9U++Gyv65rE4HFX82hbR5HFO/OhzxRZD5l2j0PtS
gIwRIlNQArD+d0VmJEDeK2t75vqh6qoH7IS/s3LvlGHqlHyyyT0dEj+clvwDqpmdcBj/kUv7L7D3
R+EIT4mhxMvJzrl7QkaDXOUANlLLfuytmU8psLusipA0UucoFRJR0KP+KK380DngI97IoPOmMBU7
zu4pZoksFqv79psIrirLtWV2uM2yu0Wo9A1NUXnLCGewaVN5cY8wy+SBWIMS/kCfn2U9H5WUttYN
0e76s5Ss05hPjtnqkntyaSsJeoMWSDqP5cWp8PONELsnKh7KxpDgXdXXCcDIk7Kw5iR///ceGY3l
j7WVE6ALM6GMAKoGVwB2Y2hRYy5s9D6PVNTtU4HZb8+jTGR1CxFdksvZ14w65XL6kVtJfS90Gknc
c6MnglFX9YEQowk28k4TazJxB+4CpjMVdbad/d6yp8FEFyANCmLgbr7MDVCQQrp80dGbPWY4ke5U
fXEO+vbkpYRXsivmkzs5407PS991UpsIkav6olfck5PMjR9sBQu+ZNrPJU8q3pMnbnwIXJYL8g1g
+cznbBQVJ0afXqQjutneePjUxEKSYVRIERWFGKGgHcpsES+YGWceh/GpCYfJReOT5uaqfgGr4bO0
nr5aJbDQmh0JNblZnX9aSlOWIIbq+MF6PzH6GiEIslW7QCJUdUk06ANGg25+ULN+cUKP7k2fLUIk
gPYzZvpYyxiJhnxhkGHMT9TzdsnCfEEP3m+VW7BxJ8IR9vDi/YluYc/YDldyj+bmTbCmBXC/D5uc
nEAQ9Fe5CpUv+4OJOKbCj8+HcQmoz/Ev6WjHIQgYoHWumtT7xIK6uAZHEN0S7iBD0J1yTrSthSr7
ZtaNfhdoNX5Ht/piLNRIst2DifHz3t3rQK9bo1YGmXNAQerM1fJd5SQUwuVfMDA2tY50YbqoSiT6
6TSBF5RYGClobXo3qU3kbU1nOJRFL/l1oTGnb7d5XJHjSxyEDhS0aFSP789s1zxjTDK7GtlkgOsC
6Gwr3M73GEVBc+JVdd3nVNJj3o9ZaTMLaiOxL9a5z4dXHc5WioTOJKySJAlx7B9mOxbPUZQaeS5+
/c55mEk9R55DzGtGfDy3iMFlm1XzsWKIoqR/ca8aTgOKiOpM3cueua7Qb2BmY1mMCVhPfeenOt5+
ySTjP/2R5/a/OjKjynNAdLEFXIB7pXYyHwIKsU/gbyRWDz+K7p3VN5XTJ7tOOvVF5N217IYz5rbQ
zBHkPbcu2zVbtasALO+/zbg5xPOnnAnimL3sIYcGieBT5UNg5CLj/yzGdzjLofNq0xRYlNaNmIb8
XbmD3JEkhBikAP9UWA3a3SSd2tU41nuoaSL1x21UVUYn7VGqp7cn3gcyTH+eq/8/JMYv2uzxElN/
SrXc0Z9aVtdtZDEt0/Q180c+07CjddbxuP/1MgfJs23vNeOwtN0wT1nzJzx+dMeFsKWT8IA+zFWy
4MzDi4Czw4yRdIeV1GximHi+gTQuuA41pNgDig+vCWbzR+6aMSU3KMeLzYFz4du87TXH0n4fYGVw
kcbX5noH7eW5IEtlvUXl/ej1fjU4kKIt+vAts/86klmypT9imNcZAI89rla47jN/YIKCeXkwxRBH
l+SYDgPE230RQtNktMZ1htAfLs6gXe32u6fMW6zyMC4oYAQ18GeEZgUc3HgryULmDtgCjs7ZIkvX
Jy3pOfMsjh9EOoZxaWfRYPwhxemAJt6vrHdRDNEUA6HS/hNJq5w3kX6YX5UbDA4LaE2oJM++ITBg
ysd6yS2B7R71Rbitk2LWTHV8gq/1UXXlE5O1C5moz7gkyzndU59Aw5IBiliTRlgYAQvvtbcUvSkQ
rbrblmrEpzeg0DEqeOT9NKbcz8lal2mc+gxxlf8G4BugcVI3/lCQfnCfLhr4CTGCC8DrYcFBiO39
p25XSMNFqBY/PLgKFL+GCigV9ZF8rTnaAISYOW2+w0JSRIXxH5JzOx4Ky4uDztPyWGVYgSq4cOOL
9MVTLTs9heGJbhRy/qtF+CpDivc7ybl64mroipjCsJlYKC7jKBK0kTCEYj9MoDBQ4KB197BVT9Ld
jyCGw8Gi9WCVE+27zU3bizT1Pnsc14oTBHP6p55G+l02CpC+yJjc+YgS+R29A5Hbos+9zsZITNV9
96jUCKcDC+uIg0FVO/QUoy0d70ldh+b0LjZ61Esk6gq83LafNr+kVP/vYBD8lJKppEVwmqMWQ7nn
x5uJ7VG4d14fF5y201UXXc+e+Iieupd/Q8hIRPgGgP19jiWIcfHJKAzw3CRwl+mVBbriIUB36soh
oyBNQMdFpxbGLgAUZBsmhUM378uBNh2CEz/WpY+ftux12tJEECvhKocP8gLY1ifWxqekmDO3Satr
+/5t8jH21LzbCRLvyMOaxuFb8GHi+7SJ47Lu+jajboqLlAPhEqrYt8wJw3bwQ7d+5OyJ2AkOjxnh
FcndCD3Nq5plb2D1AERkbIVsBP/gdVS8rfoM/qp2Mb1yQqiUyFKuTbL7NcUacnW5B54dYbwQRb4Z
O2tFez9E3AspT7Q/g2o5iRKjjZs4BO2VKRMnhPhoqhR07etKezNXzpodDOcX3T/zWrqcbg4nOw2E
eTY1sojspo4fVpXTsMtstcJEC6KUseFir0oupaSw/YlJTForUepm2o4H3xRsY+tRkkb3JFYQSvsL
kqg3BGjkE+SDlJQ8ZVw1XN7HiiSRIhnoiXIp5lCQmJqRuE+gT77CpJHAmerZwnK8xj7LNzZTvX8d
Dm+tRMgO+Zo1q+vo73AyaMxPWc/mtcY/ZpNEDJxxqxZAOSogANQ4Ev42I/U8WUK03P8Ns2EBUGxY
qfXOyB7VG5kMpQo8GSFPcLeZmi7MtTJKi/VThVAvluqJIwdnrNzyRIXnltRd9HyoRnXPh2RvJYHX
H0oyE88sFUCo1gXB/f9qkhiauR1bva6Uht7PonD6y453aQzMwg420BpnL89ANkdVUUDVZO6VpaJf
xXDLnmPUHdHqIAOsbQjxFPLIaNWslNn12PQfBLKJPO5V0pzGm4W7IVst5lSEqfFlN48LbWaKCKeo
HB2Gc7rvIElURUVlOkDgyo/kWFqclcFl3Pqfz+47baOzADcld+EJzJd+n2+/BaFMKpx6XUbuS4G3
IYK5lvdqpcB0DFbJCLMoEtdGmp/guWfqnOnYRH3V386oFel+IyTDdz4+2hAcZQORW2dPETGSjREH
HkC247fHinV13KFRlU7Rslv+rx42j/ugIMCv/jBp1jVsqP27S+KbuoeSRv9Qo1nEqTYcZQ7Bw+EZ
cWraEuwBebFJatr7qOfZHbcjPHVdBh4JOGY+XfpE34GmGWtwAu4CgR3ozCbi6kB+EpTrneAjaPWC
2KPJiYgWzmgznyw+4Tdu5hJyHsV0jZBymTHdX/slUI4X+FIYnMal1Jj6Zlh49+YJg8BucG2da5f/
8hoNZoY8cjJasoCV5ULRw5ZM0eoQXbTsAfVb0XO6ls8pu3M8AnTYdYZpmPM4r0JpsdSG7boEl/px
xd8BW8Idc6TiB4neq63pjvtIaytg0Uipdgf3H18hePsFvCn25AvqYdooEm9DXYGbrsCfN+YfB9vb
Q0DSMPOge7FLFP6XLVxnKB2FXFkAv9So7a2l18vsMLETEbafm4rV2IFiZYmZNVJk+SR3LWX4ItsE
kpHsD6rIT8MbnLpobD7wVMEbVopjU0geWGGZD66fvMrbBsGK4sAf+qh7PTrNxnxkLokN8dHWPGyi
amA5g6+EppK2LRVwxMalm6aDfb3Rkr45W4O56oVnBKPgbPEmXo1nGU5WKN+5z2CPk8iX/HK+C2fL
1SE5tpyhltIvTwiTXGrY+hPodMnlCT6ZsBPFXmpFyf8dw/bHYf4bvVZVr3aI10wrf/Fc2kD8t5cb
Smuk9oqO04PdaHxp64nB1jycMonICja4oSfrVZLpmloKyCkWdjgv13woX+AV7TdGImu5KIbMrB31
1TxNVPnMVemT3ML0kkokSe98+P99osisE5lHKqTv5OjVxYq4fteyf/K0D5t0Ghm48HyjwMCxCXw8
19TnH27Wmwt5EHORuFVyL53m/rgpFWf/zqU7HzCVizLfN1+dZzA/CJ9cy9zNV2GSj8BFEPKkZEGW
5qDfx+TEqM0My0wC5aHEHLrqSyLERXKoTnoXuoCW2OcWVsV7G4ZF0Jfv242H6bixcGC13j3IPali
Ww1+pYxY/24XrXZUajyJCY56P4iaA+VwiMYpRzboQQ373w+FraGnb749ojuOwOqQr9VN0quz2s88
osTcRNqTAk5M1EppQ6GAr+xCMTRz1r9Zk9KFmBws9fJ/Q9LgyJqLGj7KKy0ZlYX9YN8vrQWj0Y9p
wVOwJChZeP15SHNz0V4QT7sAEI4oC0mpVouerMOxOrBTfuxI1XbVyJBVN5mvQGALYGeBRAkylXe5
R6OKtG1ulRnSCAIB6uxmzUHhwDcMJlSnyL0mW7jmKIYQLUrQbiVrvP28dybhyRByZ3kfeR/NEMqE
pavEor+F4YDpsvMcNf1GBJdn1gDRAKVvkWaxV+qX3snwx3zw1bZZnwkdzQCxSYCvpdlKnE+4Kbdu
X2wTTABuToK110HdIRSg7nhL/8pYpO9p/y8nvvqSciwHLDi18iHQUReKb8KUdrJR5uwjz+hLFuF3
6UHBgZrzWvNwmJbjIXIo+3ww4n5yYGlah4DueC07uqcWu4ZH0fU0+CihnLngRwkQE89U0Zy96Ldl
hP75NqPlCMPpYi5p325ya3NvJB3OcGOk7GTJLfyB32IDpuAEFyRaKte6/A1wKia8B7lYIwEblvv+
FVOVr7KTHj82oMOIvqt8qMMT7pvCwkxm2BfSpJ6R8xcCLbKoUUXBdlpX9tOvwvDHBAmCU0eKkYrV
CZA1CXuGa3D+nUCoZWcS+FcBcOI1y251FCcNVMR66Zq+LN8q0SHegfFO52e/k+0fVWlV+AsOJTcl
wVOYhjzjkGbt8pSYzOUT3YtMPBQ80+zSGpBzOsLXl+s3ogzKU0mNlLN0FDkdbJ/UKdxQirDhWN/h
8U3yUdMhRmr8H5i37DaLsx3kB4kqF041VLkbUkzjWPQi7dA/FCKbdGHC83pNj4S56OE172dhYTCx
XfX8A+Tf9y6/2LoxoSSN3fm6Gk4xsiqgPl9isZri07kqt/Yk5gsQvLEVxSxoygHzTtRDsF9a2QrH
8ZwlFhgzedUOYYLcaNE87hNIg4Rsm2so8fWfjfaxgoOoQKiAcs1nCuKLeoDV3OPc5Tlof9fIWLvm
eKGIMz5CXZUSlyAdylKIpgpvji9fEzSKJiO2bYFr0IPGAC5+VUinIQ0crbibDN6CCyIkRgP315AB
xcPK7u86TcoVk15LIyfjHkSmNgZ118T0jmB7VwEVpXTuyI3TuaZp5Pt4R7Qy/ejEGz+rU8MXzvk8
kqMdVrzGvqI445eEV3HZzvdemb2065kr2zSuSa1ASDNfexZ07kOYVSPJqcORXmrbJYP6JdnqE3Cy
Km+QhR4JB0bdwohvwT2w1ABK+ZrBBoXhQZlp4UnByyq6ho2qGU8Nw2lUjim0pOjPaK5SCTKocDq6
NUTSt+YwL2d+B0rQr/Psq2LQCFc7w2E9KyQbFOf/dab5K6HSALL1eBoegUR78euNruwtw4ndmVaX
EqTTHa8LC6sfaCpUxpjzr1lqHD8z3s7znCqRHhlH9S8O/j8W6E78jSXQmWhr9NmuvElDYum3AiwN
prnNWIuwEwX/zFskxYopJI/WyeppvVbMYv9ph4L3urbnxKDJFINLZyRDeQOMLD+KPpz01ylwm4ak
JCiLaClirco29WZ46Xe8frTAbR411uL9AvKEe2TJjnrJcgNbty0M2U61J7IxEE5r7id7T17+GLf6
Xy7rWQ3//ePZg6gMXvSaDyoWhy5qqhU/uX2WUsM01KhxxqhVRFkZMuus6OmTDrpYc8YPqKOk5k0N
k/Efe4ZCIesDeFm6nk+sjIyZTj5QNZ5qtWBLpksnhYZ32LW95DzB5EnKlIWzQpHERfg0qMsWBFHa
4wueJIVn1LkK4gSJAwnjB31t4B8DHtc3bHVKR2KiLyQxT1OSG7wFAuNlE8jVqBzv5KOLdkyIrssm
yFoMwBHn5QlGTxhIsFCpvoufu+15THuGEzQEbV5oRi2WbHqzJp2iiFau/uNMyHef60EATtUU8Q23
hzG1qmW9DrLYphD+8oRMXGEvRNWL3zNwILFqA+X9g6zWNb4Yim2TAHnOpEAyIsGUdZKfYspbsjZV
o/gkTRxaJkwZJ4q8tIlqHvFJ8p7WG0LSeK5jcD06StvmLIF1eGDeGJxbf3zWe9ifZfOXenwTcn9t
l4OngCUjUhyG/4k+BVREjwVpKKG+c9+01jc27y+kJyQQ6DUdvEXU3QjDWCvmgU6O4VU2vf6uQJRb
MDLHEo9clxuH7FBgB3wowhJY8eDSdjUY73Cab7PGbxwUdlh/1txQ+o5HKxt9VIa01C4liMg5RNgh
90Q7XTOQcRFDQTrEZAmJH+TBUHOXSz6OduaI0Zc1165MJPxsaMZdvDv2f8Jt0zZ9Ci58KdmBMMB6
HNOTGeUvrK/rQiK1HOxoNYQJehMYtXxSnurm7dBJhF3NpTD9xBILGKby1HkbwM3faUQ+4H7ki077
BE7HRKK/WcPl5goW8duH7z0tROODTIJNYaGCSE9wdQW8yGB2zSniNXzv0SC5w+82u7cT9L0ubbuA
hKcBrFVjlLCGllRS5Evryq1sywhFYRkVKTqiZ61iVPSH3Z+Rwim2RHPLXbQyg9cluPVmUsFMd4ds
tJOOWVRnFsa/foseALInrgGYE2EGdsJuRJ5p79ZuzpIw5fhuLKBiSOH7ViThTsQoGRzsyjpxLrj4
o4BpEABn31955lyXV9aNeWvvgOwWMIZXEVffVp/F3+MCPLTlkpesZEGUzZ6NZPQTevaH49qbgQ3W
59i3R+fKxzlUsejbMCtXXrqxvav0u/gl/FnGNuFeI5tHN+ikLwHPkjMvwaiYd/dF5xEVaE06E3a6
aLCLOZZj3y4kXV9Crq97PegoALsHnlYCvn1vEWbBhQXHcKTbN6XwSBh6wR7zLG3os7/LIyU9qBzc
fTrumceugEpcVCQ9bnekbZCDKwdidEmlEAOOPs0eIvkjH/j53kbjwDfXinvFxdEDPeb3uKf0kLqj
8eBwS3wUggsUJ9YRklFDJjVMDxjOGq6VNLIpQwOZxgpnxELnKrPVHYNc/vBhbJh3MJeogjYJwNaR
STBjGd8wGBOCuXwo0R4CWSj61Z2dSwgag12iUTQUiy782gFt89RINeqOHfFgAq1vkN5FKQTJQGfk
1e+KSOTjzshC+MAxIlyvPxrHGhQ+HaiSw6Dog9BsGSc0DQac4Di7X/tBkoH1NxvBzfP1yVp1ivoN
vHspeu68mL5U5HepSMBN+L1p6f1ASq8jDfLSJfuX3FbzseC7A7QJ0CeHmy6WRsWkVLz/ij1cCx+f
sPpW6/iHA256c4p2XI9sOFN1T9lVt4xTpwmOOO+s6m82uKBLSzX09JOtLR8PPrZMRJ30lqgy6fWc
MA5pZ/OpvGbxWubIh8bpNcIEczXEonyCcW0B5Fam9g76fJMRZkCvCig22QS6AD3mYwHV2vMV1gmt
0b73zIy4S4MXstXQ+xsScJKfaNNivmjmVADXcLCzzT6mr6VqS/zQPhh8UyXxHuKeGmNsEvY0wa6+
77A8NtPXUuF7alYvLIE0EkB2TzoYqoimhuSPVCvBd7fIXZfXxXmyRj3ojx047wt6hAC4q9sQ7rTP
UKh8o921A803km4x9HED4Y6yBhmjmm4uUVHWUrlORhFpXr8hH79b5o9kxpDJUQbHrEs5YKX8bfPN
myUXEdLzc+zlroMhrHtPdUkuZ+utbJF7eVu2wpzYFJNn6gqAKkUaWbdY+sYQ8d/e+zVK+v6g1MA2
VQnKo80pTsEfGhsfPMVdGpLsL6uwSn5mQMs3lXn9sJZE7sdbJjtbDursmyhJCLbGqsbZjhQNEZUT
QApxffT4hHRkQR52SY7fWCaTap0paVAcMt+iuic0laI7XTdOKAirI5Ex3SUCIEDQVzKVXAirb9CD
DPQGSo7sy50Adyb1BPCPpJMFCzJ5P3sapvg+cxCWjqzPxZ/kMIKow1we839uH2hwdRsABEI86Zk8
8teweFwOpW/ZRF2mTt34qC7txe5k4Yd6qe65tWO3eM05Lli6T2FVF+zhWzwqMU1jzujFbexrc1Hi
PNyhY4PzLpQDBG6ndPafpUW+NSJ/gwPmND8iHiQMTf2+ptxvLB3ParNlASXj/2qBDsFlNETVLAIp
jQ94OQ0baqtJyaCQe4q63Vzr4rEoCBDKTxZiRPWk4oZS229wGFTF2nQN8C882/GXuRN6LxfGgBsj
BFEYScE7bRKprOkD5CwygADuZGXxrEXtSq88PsVjY+nrjlqI+6UPSrKz7YbUJLA22gFvTO2cXgC6
aqd5vzjRqrjrZQz7eSHdwbi3Pe3KYL6xhX1dqHUrLGlIB4QraLvv+jsG+5Vcj16J9TseWRuRDgkV
hXHFKgjIUKBHDXffWTVL7CJlF4DJHIJIB6jgB6sPNLMXzC+QteB3uyPRmf/UjsX262FrznPEmJUF
eSnEBQgNIC0SL+eD8Z0WKQ5K7vNtbAqzqn/DR08p/BawFMmLXA/ogiV1NLQfOqubMR3nbPKrpdW1
/TbyUviP8pR5tuAEIq64lDhvFlau6fJTb4L1w6gYA2zPBoO+FtICPCYq+lgoftrsi61toZgpDlVj
DHX27lCId4N2+qJT9m5gWGG6UApbRrrM2OFlyO3PAFUa5+cRbPuHAkRm1XbtDNxM3VyZmGvp/Hmu
kx4rHm3eXGV3XL5naQvlHBiRaz2dqUgdKmxuTWw5JbEgMOe6bN2F8RAswNfKpkYrCSysuwC0d43i
k7/E9H9OEW87pSe6ErjQdQmsyvhbA/Zn3ADI+8qTEylj6ZhqpgvmGuvEL/USDN7PBdRLmSNUbYom
B/RwqZ4Kh9B5CS1dLIYi38GwMwV8Blf4H7kCLrmsEwhaCZlQGMJTjCLAHjLy/isLyFBSqHGKo4vl
sskFaIwfopRD9//WcNMJAgQ8qZtNAF+nlJJ3sxOUc7g1AO7dKBJvSYC+FBiP9n6TWcT8w+7DuYQA
Sh9O+Boq040QYO8MuZvuhKYaxs0fu/t/ZGKJYPP9tPXtLbJnFAB2DQSMgRwAEjaObGqnVTgm0+xB
GTyT5xrHC4I9o9HnVpb3piQSDD59iv89ELonbllbbjnai+EKd2LIsrW5qe0m6JNKYmQ60Brq6wFg
0K+gv6kKWcFu1FxQ9B2EekziQV5LvDoe7XTsn9UITnbgC4mJKTAjpFMRw9LmYsodLTDjsUMGXdAP
Kxf83Fj40yOlY0vz/TQ/R/7H+d7GzKp/sYw3i+IsEyg4jXkSsEW0fhAluozUZTgJWDZbi1x//Tm8
L+/37fORbflahDxQUkvl+fP0jTINaua8FvJXxfaspfZkkyVBP9iLGYvNpzeRdBlAOonz+zXo7soD
2oc5KaOVlOS6y92kZjjJcVySbY+/npI2tMo0CRqYmkcbuefPqQZsa6hgfd2BoIYMVAzH6XQxsG0b
2KicAVTTMyUXI0bJ7wuI4nKnRx1u9xPba0tw8IInBDjKfWUsuSsGbPn5XXcFNq+2lVUuaGxXtPgP
aBdvk/G9NxknltDMCC1u3sFOji3iarLrE7XNM9o8/0OZtBXAuRufxebbMkFAkaQJyUQZK6Sm1f1M
Y90lAnPZ9Xv34td81tlB60sfwY5UithIKMjReBeKR67wimhJRopH1rpksY8rJuxDUuPeRlp+pwrL
BGEiA/LAet86eiHwx38gvWqtT1iI8QqwUKSkOB4PavRjRFqGAUlgiBhcjqMsHiM4anAJwMUC5Fme
S4HbSo5BQbVGCvZLR2Jun2krmKhRERJSngoGOvXw4gMONKM989CGthUkLeXb1BlDYONpHWKV/tiE
8dckHnOGUIMTgF6blFi/fG0i+9fJiG1faT/kczUvpXX4Pb5M2PckmrTbN2JVREA09LyAEVXImyC6
UDqbOW/r+UPLwTayYa2/70+N+HBvKQIucM/AnGmls7hNcCSpCkFfMbbTekJGef9nAxFoxGZUKSKA
y39ph6KhHCWeAEiB7jGSAoCvgi1d7dpAGJUqBpLJ8kS7yrfyI3edeK4EXf4dI8KjNwj+9yrgkuat
ZgRN9/nfhegz3YVrZnYpXrXx6K3sq/GeYcwELB7qz6pjQ4U1FZDoZeW4DbpB2ZXJx8YBWKfarEp+
UuYHK8w8+1TKMSUmcinBFyjOeA7BZKm4KECwBdkNuHUOrIGFJtjf2NR1CI3ILA7oBF4VRJGwzLI/
jgHotmAWQ4nc3Rx0hH+z9ZYwqKW2ZAQmVp8zcAIylWh6Dxn1HRFwFK9+FBp6Q0STgNE//F7lzuYg
dQuTBHk4CRSVLureak/wTObTSFSKYNuZiqUQe6b3tiFoth+Nr+EKWcX4fh7javhZ5VUY0dWCGzMR
XLLhxf7xf9eA8h38kKf391oeSnjFFSUTiDe9+1FJpd7skhai6oinsP9gK6cudFcu9Ap1crCT65Fd
dUZw4KP4SZLevTX2WlhaqOAlwiQqnmr2QgRCtSAo20q+LabLSL+nSsG5Gd6ZvRo1cUs/ehJGiS2i
K1bDeMevzYcuK0dAsSaGVyM7gXpYfJrK1ITbeg2YUqas7JUymByZWGLNEixHvvfe+M/jgFAVoH8r
/SpKG4bq28ahPZnNPFAwCHHsA1frMABSOecK7luALiNkkHIGGStnR+HG7Otk0/5qiyKoOAvevMId
wMFgq7Tl1J1lzPTcqCgVN5kOUwmGoq7vkZspG2II+zRVynNqXN5iDyMlF+7rne86KvffaJsHXhoh
iof2ttMDfFsFEOvvd4jiIrZwhKf1eIq40MhkPSi7mvGwfNJmDWIGWf5i9QI8DfRZDApBK1VHej4Y
jdIiPIsWR7K0VC/uU3Zfw3Gd0+NSP/UtQBQaY2GU7+uM1lMaN1qizwvfsEhYwmvUWzTII5ov2duP
z7XeM+lctrpI3ufp14GXVXvZixgXTC5im2ZUE5D7c8BsAn40nWIlb40pUTNkcK20kJrFq1DPipEI
iEcSS6Q84THbSmb4JiiPwhqY9mY3MU/gaxT6hXIvxBex6iRrOBwtsCQmDa5d6Zy9+GhMII9LFlWr
haDhAll/xHV8YtkCGJuRt1VnVQosIwqMqweSATnpgGdS8vXGNn3LnLN7KBbTGQnGjkn/HuE4+7fj
H3V2NizePQ8DoiCnqrkf+xkh2mum1eYcN8sxaBUCEnsvJUj+/MJdJYo5hgQg/OJ0VuaEHpX1TIlO
FnLNCovTSXtbe25wHm1jtUAJfyH3zmhkENHPDTZnaeY64ayJo3R1IWaTzxFzco2uGBZ0M2fDUdto
QsFxvi4UT3AC3FrnowN3D2jMrCPPERWSoAV16ZZ0XUg1K1t1f9tCHz7z4tq4DGdjGfG16JSwQVjf
8mVKCn0CoE+btUJNFenGVM++ua7xfxMzFySUesOavJHw7z8KfcNkrmDTC6cg9+YTs9GvLrn2pqz6
D8OqDAquhKvlh9ap+E+8De8LCxp6H4aEAJ+LuCo2H1POErRSdSPOkFxwJWpL5OM2mBl9l/fUdk1T
BYTkrVHepk7Zs/CuZCOLLyh6D7p056xrDHaUWQAprLgdWqVH5E9D4dm6y1y7Dyvw6jAP6R5kNR4B
091LFxRWJjm69wvzXLUO996bcDYrRyjtRSIrbmgvqJaTbwBMBYhW6SPmo/AznHW6r38OBlBJTcyW
6rHA/U8c3JAtS/LjbKB+lk8BXPklk5aCi2ulFycQ3APYzo79Ef3YYX76eYA30+Uxk/qWBe2kpCkA
lWJjZ8icDbXSZzzrDR3ZDUCu1ly/j7b487fVgdTrl+u3Jwf+cVQZmSZzvXYCtSAUcflBiXRokNFm
esuyktazaw+DeEkTQ1APOXRC+80zKVYC5X3d8iVtMwbDYXwuzZoS5C+apfR/R8pBxQc585ydFIUf
mMT49aSvMFUgBieLW+ni6jFlEyI74k31BGOyjxhquw7aapM0RpwHxVCNLH7ueQOW92QJRqq+VNL3
3/CuDtKp1IJeTQMCXN9Ag6E/b4DTIuX/IhESCW96tyuYRZVshLJdvQkc258UzFzelZkPY1QVFAVe
DFiUaT+sW93L/AB0srClCsxoQFv+FlzlRB5PC1eJwkUBAALmYkhgjgiKdQktPU271GEFRjXqFkTF
EUWKV4pWjgd5O/PmX97niLmq8xPnnQGQE/1f3y5ERQFC1oApq9CAX+B9zXJUnhf1vLo588wvyThT
E35B2m8zjpa7HoFkvrU6PpOAVgcrwgFOvHFVZEtxka97uDSgtpVp7kLs11oVo2MakGN7EtYM+Eb9
e1hMlZhRIg6vGr/GqGImcFdPsJFM5SKvlGSMqGvRyq60g0epSaaSQdmhYTGazloQ99KU7qSzyQM8
dGslBiSneQ/0Pl91kzkbN4jOUP2XWi4ig0pb//5SezZuGetw2rikflH+4Q+0EZDhoFLTY2KR0bMd
REg1uJnPYnNYK7HzMR97/w05QQ7IYnzYdUolQUFJYaSAIAnzBoz5zKMR3ywaax78AdvqwpvrGzdx
nymdognuK/2SZJSHZmk2ENH+n2ZZn8VCDbUgafWBIOSuLwwkP2nI0cbZ7rnyAsM5sZswvE8eB15V
nf+3qkdnijnucPl42ydrHohRC/83blEo/HSfGuLq5mXJY2yi2ZSHHWIWIW1qBIfFU2KDjJ5KOYKA
3jFzQzJdhF+pvzMJQ53NR2wlJz7gmacEnHc+VmkQJACezTaKugnkWQRCmLyV6XoDwUqpJvh7Slls
Xl4CFb00EwE5atTRYJe/v3U3AJqMqBr0UKzxSLl0olIDvI3Y+m0zlqlfHq/sGCWjTBuVuxhxmmXi
qAWa9ce+Zr0WJTTP5WKIUT4qbTZr5LWTBg818mosLneQUMSzx3oUHjRoCB1Cp9LiQdNcAtVmgqCp
q6TMz/9fFpKYFnFWtDKYNrIJB5LiZJOacS6d14wo/7ikgmr1S+gYzBpHsUAGLPk8BuncYCZPbek3
pG1EXRBpR1sJQYKmmqcfc9akE+ItqfsTiAhaNemyKfIyAO4B7Q9r1gWGnobpuz+Tatg0cnTdnU58
ODdvRrr2C4S+hGsfCUgAHl5efKpuaS0jYC+VUjcT1FHnEgpH793aYVpIv4QBiuMajFbBcWy/7Uvg
Q666cNjk25Hklz+ZzbdmsixeaGzZl6DRWclQW32Bztx97NE/TYoo/3kRo06IvkvBvjVpqbi9a+aH
ZeN145ypgaM/x5r/BA1U3E56O1p0l8kyei6QgCa4P/ueizmXRDjK6o4UtP+QHFwzsLBV4z9uX0Lg
lvFdgpVPXIMo8ikDiH2lx90r4LDQdUocfCILDjiAOT2f9uu7yJfCwvbRgUd0dvAILXhP+/o8licd
8IEXvVzUmpcag43OZ69hwEaLD5rKJ4TnVgSExtX3cP1wzFZTXXk2TyBRibKbL5mwKJwYdkau+4vH
yaESKw6+LlnQBr0IB3rszSRzyg+9lgDJeB8q2cl8VBb0Kv303tTduPpY/cep4F/TxDtgR248AEsP
Kmb6xxt7lwopon9u7E3SnXJorwcrV9eHQ0PgB3GC7s5KfUGRDvvfjc3KMZkEb3cjSpdqVFn7z6Rt
jVjKyKxvZReu0PuM76ZiSwv9X1093RLzgNDXe4IMMIGAE7jSFjQo18F1gkRv2Hl6QoLwCr0Ktsqy
Y2Lx3PCy4YVx/NbhDgMtS6GqyF7tUJrtKRHIbIXNVUGr2C7PokO3RPeHFbRhXrsr249hPy1dcDbX
T/HqwARNAoJ5wF1SQvwGnEhNnx2XNTGCKzJBX3YntztEDgSQfh0tQNDk5OQi1F5mpOnJM0uNR8h8
8nNav+fLSdfwMG/81/E/Pg4/Mkt8aAH0b/XhYgSXKrFwae4w4CUziBRVCa+rPEYjBfj8tW8Y2VUt
AdYAAAziYRRZXRlwb3+txShDk/Jzrg1oeodepa6QLsZ3VuEE5/4uPkgEB1zNprUgSUeE6K7aXKmJ
GZXvbH11SLkAfoaYYkNN4Sb21BQaTjEGwezwtwbSxuOHTDej0Z0t6Q3WCZcAGNmNX4ZRS+swlQrm
iTlvh0I7m2DGtRIkQZusLJ84ELfXLcD9BwMzRlQwzT7OR4XB3Zsryt003LJpXIEGhxb+NSgVavrL
Ciw64TAWWx4qCdMk6FU97lwzEgLFIpe7oCcWFTc2CDIO3CNXs1etH+8xuM4x1OVVXaCMqjM7EhgM
1HVc26+UX9D4gM/l0/QWoV+aeHe4WmUI+tXyu4rP/xsx4lNIaed1Rwhoe8BecikinJ5p++sSz/AS
WsVGJAxrLxeah4PrHZWh6rQP/fsWOd/ccM0zcjnlDz3KEP3Hft4BVoDRj+S064z4d4qcb8I/yHpG
R7kosp4UESIF9e7vx+ld+iKfRp7mswGwBvT9PFxsQ60n0bI9tZx0Jzc3bhqyVM8Afi0xCe0T9bJ2
MoT0Q74tk4DuA2ZzLrisaqpM00cYVflG3d0vp/A9USoj22pjcjahw7HWW8cbSdFUHjmfmCPS9Udg
R7BS39kiBo9UiihAEBMr2PFqqM1SWV7xwy16SMIjvj1OFjcTMMh5xgcZuf4ixFP4Tzb8blfm7Bum
ToNvJHy0AGMX9iAfNkGIXhqCP2v4ntIfMIoSSKFad9ukNgKmVj6cJ4e69CFLIZyhUyen77ZkHkX2
Hzk5Pm+7fNv+N2MiypnXy66PddWeYfAfX8VQgrxhChtzQtZGH+EmNA3RnbqZXvF1AIYetJyhZ7P1
fjDca289nX1NfU7YbReIEJfEYt9Mq6hWU+GW3mTboZhJzNyDYdKBbKkClQ5N2sa7TrdRQyxAUhsU
uP0pj5lmUc+KHwMvowIKxCigcHnmy9HcqJC/oQ3H1kl1fi3PgWyxDNpoTBNbCbWx9vKwfLbE6fH+
hoBCIkjzqOrUkDdwjxAiM72xJntCRM+v5kHYurANDfZhDfHeEM8SMCPTHdCsSQdX7vyILaUiP1U8
lNAU6iw6Ha+v9jHImWYc0UQX8lzis38xsD7cjUI4FsMNuucfIpY5IBuFgMy1YIgh4GDkNbpmVCTX
PcRUcQEcR9l1TrTwAj9GlSJX8GpOkJJB1PzTsF2tEKGM9iaI9hcGbSYk/L33G7wtmJtzBa8h/pvg
YaQSO46aajvU+1nern4K3P9x+VLr0E4KFX6227+2YU2Sdy6dGKpTHuYzEJ5fvtm7jtolcJbUd/I9
KQEOxpmflNCZ7RCY8Uxlr8Nsp82pLwC67QcfNyKf/5UtYUvDhRQiTqVJ4IpNWLIEZePgs4XA6tIm
4vp+UYPkNWRfuXkioeLb2S38ETuVlaFkHfnKaJFlhZ2hHO8zm3DneRPraugcN5ibu360wtbH5lPN
p8Xo0oys28gGPueGDgI74d5w/naaBefY+/eYMKnTIl3Z1M8wpqikCuG8dUhVuWswecXBMae3DJ9H
qUtig0TzEvWIHc1xE6HZCyG1OJwgXWc5AkQRpX79IktNyfSPCz9iRe4uPB3jONUMdo4kEHTmCS+U
ayDA9C25+K3tTvBj+96XoKWMNQ6vCqsgxLKo6bPWOakQz2DY213li+sE83T+h2kO9f16+88qs//w
8FvzsZukwrGZwBn4xFMCN6LuZ6vig5XzOFNgc8hxtd1e2NazpGxViwnVN0TGJywsW1P9ziDjSSRg
WNtdjsGjyECKiVZzMGNFUsavOFyGA7Hivz5S5DLcptnLTD6sLWT2cIiqQQ7h+Y00W567TqH+32K2
MsQ2nVKJi1+urMiUNyH/KRz9kFSQYXQ2ItyYgF02al+246pEKRKy0UozpX4qvbRI5ZT4DaYwVhFP
5Br/jiUTVwSP4IikHpXbNnxzd/SX4WOmBeCyPoosxNNHuO1A+Yd+x9AiQKn0nfNXb0esfZ7gqaRQ
K8jSFur0IeyakD9Na+mqJxZKA25h2UxrngGlrYxHcmSK33z4VCwaRRSjlALqDqGclZha3ci0pEdX
QdChIglUVvYJ8AAtscWwqlT50fDX3wU5vJyT1D+faKLTSrYuUfj5U4V0wPxHkIV5JYar34kDCxPf
/cfRtjdNHQeUzxjjNt/dcNzhCBw03deF66x+5TFgihmEINTaz50mSHDWG0aSuk4XEi+Upqkw7+Sl
pVdf1fcpGkOJuUaHivKmWGZ6DdfSNfvyE7MTgy4wirs3b9W+bS207oAAQra/3Lcw6cjyY2KDu0j+
iOJefVvtIsmKfegkaPh1hFPhQU1rHh6Hof/8k/j45Nqa31VymTlmaDcL0k6TEWMkPi8mWsH9rE4H
F4rJ8w2uQO0bA4JwhS+xc7l0Fm5F/R8BO5m5GXagrBMUFqNHyS+ZHg5wDljiZ0l3Wzmpq1oaqYAb
cQ0JGf/ojrcSWlp1fSdtzrBlhpyhRWnBbAkmfnCcAdD41l1on0cjmD2Ay0ttpj4ZySQy0qc/qXJ6
OsgXH0IfGLl+V7RG1tM9eduOKaoAwAfH3HsMbe5J8qD/hGT9iZYhGtvC6E5AlCCNwNg+STWSZ7vr
NJkvV2Ud4TXS5/Mklrkp/zAgEr8GlTBJOoMN7tbhkonsOVwUzvXlTsknTsOSTfjI6YvOZDU28Oym
y1gIjiGm4qIMmC/+2DSC9AIAtNFcZBVTaJmP2huJAxd9J6y7lUOpSbWnQnhGED8OY8PUjdsKxM6t
9PEOatyRb9LFM4VygfnCuPdhPsEo9/r3T1IRMhJjNR177f7yX7ArQFqTCdYK8qgy1hN/+KlQAjlW
mkFLewiOVkGgXsTGszsle5ITi0CWWZCTtjVvZcYiC+YFyKjEMFfk0qZ1x1m7ZeWxwa8KNVnQIeZO
t5Lf9SXoOnVbGdkXjv1S2hHlQttjQyjuEUwZVs9Z5o0HwaJTEc2i3b2oukEfnpwF8v54hv5CeO63
SY/a4+FUfQmej79Gd20NJRQC2+fevbiQgaUoVECfR9/ybDKgvcT9vdnAgr13kpIxEGX9rIKoFxVH
DROLhkMS6zQD+cv50ijkXB7h0rRY7uyo4b5iWbMqcMbZT9qA5Wp+bMf0M9mqjEFlr0PnOqiciz+A
wx5MDNOEoeGMvuIcmk5zWfl0SUJ6o/6XYTZhMR8ed/VaQ2iEieKX73c1Bpn60o0M5f8YflmqwH9V
2NN9ngvy1j0Dw6umybLQrsIE5wt6pSnKigWJ2l4aFXz3bTkgm5d8hKpm0ouhq2lK9lWUK8qiLp3T
F/tTmZxyDsE/os4HJ0HhtYS4iUg3p3rhCupIs0sq+HrBrNfijTbiWQZ10zZe8km8VHtHJ0TBeqtN
xTxa5Cf7SUBYZtKbSYZ0v1dVCyI9jKB0aMETsED3oe/8XdOBA+ggPThZDVa/vNPSpNVTaC1NRsuR
I1CUXoHzmk5Ag09U21VXMYdvOI7q68RgJ5l5aIdCvgGvFENi9EvZ6NeoxdPNYwVtK2XgmxDwoaPf
PjcVmVY1b90MPxo9a225eh2Q/QVKEdxHPWtUihjvrd/tjW0p1AV+yPUQcAO79I6ixUwPNv+nTmtl
MC0Gktq3EL7EKAilFQ3zZoRlsch4r//a8XnVOLk2ejQwVwg+u0yEW9gEhjpZe3iTdSG8ACvsgkT6
a+B1vifg8IC61Vrl4+2zwOYql6OvS0plnD5ZWnueE28ClWLn7hu7CR1HD7DI2V/ON7P/BYlgyzfN
G+5Xi7awiCHMdkGSwM6F+6wGSC2LA6uBXsketSWFmIgOKQNQy10oTzctvF7VJOdu7ZO0oA9NPB1+
CTHvwXWBNN/ZZcY8Hgr9UeOZ4LYFglvGepe4/rYvwLiTw5SmFJWJNGiGDEOj8WhjGt03U1n7KtJF
7WDf65yXeCWGJcOh7KWrXk/QMWYM0jixwLwsXM7b2DvyzpiSkBGJTC9QuuiVwvuxVn/Yztd/6qcP
ReaIERhdwuwoo2ys2nqtIJinUogdbFsB4QUXWWnOYJB5fMoao15lz1dbC5EHmolbsPJRjy1buuSC
LsPxPftnzHS2XU1uI2BOufvDm9wIBxb/fhGKqCahkOXqvdZSgLfzRPvVTCmhF8PD23ukMaoqLxaJ
pIyNkA==
`protect end_protected
