`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Y65/MFXWhhADwOVv/M4+o8eaVO22scaJrgCxDXOByJVk85241NyhfA5m0IyE4wQJmggZhYij4hhT
+3kX1z/WLw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZkenUivUwQ4WI4NH09hs8kGW6MMq4uVGfw/NDOOC+R14rbma7ZeAsZ3KqSxlJgje8I/XUuGZog+Q
BqQgUXa+ZgnYgmCAp0+g5H/YK8jcG2T9DuF4eM1S2TWLZfAaJ6+Oih5mPKEgnSN33pe2nuPG/tCZ
WXp1OZFZ+RB/28BEUq0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KfYMeFs5V78k6nww/KOz0zj+63zNb4UOtAYickTFxZ+X2Bnwv4bsMA1cXnQyk4SRjC7e1wBUUIR4
UfTpnVYzTQ8JpcBUueX6sU4fNn+O7u+hXQUfZAI3YMihyTW0Qh5TEK+Y0Uey1NL7nPsKoI1AWQ70
umGRh89sWKiT/oKyLtcRew/ZbNUPpJUMKp9lrijWopqWCeA5ZLFHUV2A31jPWLd6eOES4Ksq6rju
hbFRC+a1t8uoCoTa2PZzl+q595bGHK6L3br1Ee+Q4vWmyblGzhWm0BAImBBFo7rXmogRR9sSFa7r
Pn0ukX6kc6eftG4ZTJ+XUDMCau0/outNM4zjsw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a1bFcIkZo4zPJvMJud4vhE1uFKNbhylkuzUR4O2EkGwLrE17fGyp+MqRG7r5NXGWXZuU9WK/9Gjk
0rdtGmDcrDBvQvdIzWLM9suFKzfFzhT8kOH8hlb3G83f3ynzmwpzUUgKGmf7tSHA7vQcdXCyq3MY
kFp+tB7AzWsmU5Ifzj0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wS7l1EcN9oGmeOh2wHa8aGY4hTUVFraqFIuVxqm0oqEK6gJ2RQD6ljT4vhdDVHw5uWV27xjMC6Nq
3j6hLI5z6lDKEjZm6dNt32pWA6dw7FadASbVwuaCyLQwHr+jXMBETZB6CFmopdxOWk0tjAmuNT8S
6rrK+f1fNYptaPKfOjH2eU7LJItbPRRhiA0sHPOwWzftgFEnTC3GPMw/GNmRFIVoNJWdXxbY2F5X
9jIl0f1Yz91j0MvUjp93SfLG+NrxinVmKZNyCPJxurpHvwOuxUesjDXLOc7aaF+A/2LfTEk2hzWV
MhiTwFpPJdDm6LIJJhpCOu3SBVA2U3JHuMoe/w==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BfNd2bDGBtVeSwbNHF20kdZMav8Ejx5EwGOiOgAGrQhSyAHpuGt/EXA501iAxaGv2XOVUgjVCInS
6ZqAXdnq8jYBca6BFfB75y3N2lAKe2aXiu1WWsOyb6BrcIyOQojTYsLNE9LwQktidMkkFBM7XJIj
HYLWwK7vKg9moWzSIe96UK+ymfjAGVJFjMRtSVMdHAbKrQWC/dZH4cYbRVC4BDkNzqV37knm0PDx
L+DaSzp61qE/otP3FteBgrxdQ1xkZWWq18DuN4gKD+tcxw79LCeiimII2/2/qAe3L7sYLPUZMih1
XflOAcTbAMQkdolvxpm7dxjneu28qIJPdA8CKQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10688)
`protect data_block
ZB9h2BkRgORVefM+y5dAkVRcVpxf7ywVfg01r8WBKBq02uTsfoRVfRwXg1Yb1Zh1r2BDIfFU5n3F
aSScauUQrjulRkPhSue2hMW1BgD9qACoD0XjVFNQOiz/DNAKRHn7TgE0UlFa+T69RskpKnjYjufR
Yzyd9YKYXqI5KjyRCkdcby1dIVZWhExV1MgNLEWFVdOf1fKsomjRxb9A8H+Do+WYo8Pncyb6PS+I
ZqR0TlOsCkM/eq4fv/MMzvq4njkUzBx5CNuoq9DIhCZfzdI+TKOVasqWUrUHXw2TPGr8OAowZZuB
zuYLeWJSYh1v+omlN8befXSDXh3S8a8QhyqsRSZ2OeTiiOdWJplGuKTUyMn7GM8MzHtYYTfrfwcp
sBc2PkCfAuq7oiFnWqJurRhOzw7t/a8L2mrXWeN/F6GFU6KDMlUqDmNRfY4k/LtBqbJYifYOtLXb
R+cb8vLj3AEFP4d+rqVHGSAOsbOferso/YzYRv1VCTbNbfCI9LIFBbY8BVEQN8Uw/QBgs1zDPxJf
vReGtir+2uHujEQqYyzAENYqDApFgy/aRlB86xOWDbocKop3NJeBTgwVBpKDucvkxdkdaTDRy16Y
cAASUb3XW5Ucff4SMgLyBmY5kH9ZYvKYCI3qgASlKm6R3RGTD1YPvreQIpuMsEhIthFV0gZ1qcXX
oat09OMJwc4ZDsa3+4G3BSW9aoM/sbQZV9JaqieZlNOAkJKKU3cG4T2H1ldbRiUUiWRGn7EoChUl
N7BPx3xPWB5eR0eK2BM3W+P6vvB3CQD8nq49nwAxwS/0sWy7gNEh/cJyBi/xTlymK1nQ6V2a1p05
Zd7eKKlXXZE18fl1BfsqtzCtKM991DjsyoWaZcI1vhGqEgKGUX4ICYBqJMhNGjHIFHKou1yCtMHH
iUyl+MtDPNOvBhVABeFfzaVxJRj6LrwanfrNdtiwG9fPc5M1cYkNwso16JY2b02qbxbAw3AIV5vE
EhmhZ+P5s9mk14XhQlEiEmRN1Pn7yFOi6BaTwE2yHPEGFDvm0wHHeC7P/bBykZsN0H1pCAG02zO0
Fl55s0vfRKY9XXnfETfLRdqs3xtIQLIvE2s9OSk/7m+EeNTsCRQoTWZcnaTCBe80A7PuIfCgmKRa
3NYLPFbvH4ON4HjbKGIzt13NXBCkpII43wEZJaTOSSnGldijgw3e+eLPpLM0f5SmXjNkj7wVjmrS
ZtVKTtlXRCw9155FpGDQFDpGt9Cq2+pgxIJACigzIIEHb3fWeYd8KavyyRFqAyKo8y9Mmxc+T9mq
7Gp9bTfRDgawbUp6+Nes36f1+GNFLohAsPABf9UnhqRGUCVeaFcnchwjNcxbi1OuKFwzaJlm1VPu
DjoRDFiewP1hOMMYyYLpRHem8UJMrRCySvSbxFjhHz4fp+6ciDSofY1IsdwsqnJKtdkoRVPP7Zr1
dS2Q5q0jipZfPwl4IOyYRUgDCeyb4Q9E7B+9M6Kwk8TWL44gdFPpdxSigcXn9EA0p2CQOO+AIfxS
WmNQMe5jfc2fbTW8FjgqipyCXVh3wYV24yW6VpAEmeZrFdtNZpyM2zcwP4UxWa2ZYMqT5EExoBFq
ocU9SWW+7KNJBrsyTkPB7uUysN5za+aUaKytvSy5zqXXRBj1FcijZFt0vzu3D5ZinRSDuYOLNE8P
X4StC32AnuNOIvomqf5BkUAfveA+vJvyb+MYdQc1idHhnfCdFkVJxpEBTi1wwA0MSXsH4P2CtLGx
Y2ReAWbwuwdhRxalYXsRGUHmgGly5UeQLkchzhlkN4QgHEGvlbBLYkbn6FmD2an3/k/nFkirNnVs
bn7hfzL6J2H1u0439BwrJpM8K/Ne1dSUboYKtIvU3+dgB6ASPF5zJElZwrcW0oTsofAinWC0ViCt
RJoK6HF+aF4q5PtYaf7l1XPFGPL5po11tGNQG79L7FsRmZhFUBpOySP2ulqM3GgBt/DeKa6RSB8p
8dbl1tDokThWjpEZ8AMxB1QBU2ul5/3guiDJyHU6gXHRmIfyWj6yEGI4AW3vATgK7hquoRc30iFI
0nQsVUFNT0GCXKrTqdDZtrDvAcZfBI+6cAhC+UbIFtGKyqick1ctKGCTGFV3O3UT/DjzKO4yrWvS
z9PTX0E24HC89o0gBLMoN7h5fneSzLW7o1+D1bH5b86HAF24df6MsivedQVzKgAPbGbRP27jNfZd
jWMlTD6s3IjpWM3gefgZ+QsRdG2HJox4S4fzr5raS4bq+5vhMqI9X205IWz96C1HRr3VVOV4WLK4
mHloBk2sOrZffLEspy45xrDk/5tOHhZcLnWmmSpeHUBZACWmWLW07MO04l32oNW7qdGPBgQ0nYDU
Milew3D+wMo2vWQbyijRLb1+izA9NCX6MMyXwF+ovnCn+i68ZUrIALRM5xGVE/f7+uVXRag6k75V
keFELiK3IrZ71IxyhUH0IA49xDCnpXj3fmaVbqTmOXSXGoRA3fmZ4nl6V520YhmEF2Ig5MslI7ww
TZzLG1zRCscNM1QzH8uddXzOr4rOC0ihOPDDxG8bJy6eO0DVnguEhIfCCFkZqb4ePJG1xwDuf7eD
LKUsyGvs/hwSYLxMkPT7x80h6K9nXxkwtPuv1DcLRcyY8XjnqSOwGHd6a2PvrIjhijKvY3D01bYW
23LK1XL6cQKx2qM6IgH45itOuVaiQaGC5S+QT7hKhsCp3obf5avgZ8vDQScVeJZz4UrwVjhau4tg
zke13vkqAb8r533bgEB4FKYSmoScpm/Qq1fB/zqz0DhOVtIPZn/F5dpTwxuBe4vlBnbeDizN4gU5
eTCasiv645He4rLRkuOCdHALnhQS7wO7ZwxNmDL9xHyF7db2JH3fLv4niL1DMnMWUFww1yr2bat8
cKzXiddFqn6Bwkb40s49LumSEeP8WDowXo1N9EwJ+SlEgFaoMsZWdBH95r7xIo/iHoIwZiskKljU
UgqzFvL7eXv+dRFkBjAy/7xf3yC74Z4MpvvhBppewzuVo1D0VyfHsNCzobZ+H7dBcU8O5Wy1SNRZ
ESXq8mqqgX5AoQbo0WBcgNhwiSSCoHiJfJdwJm/oJhFmNmg2vzKq5c7KtX7b1S87umOsnxDOw+w+
lU5bzjP2LPdIVqnq1upQiD8zlLoy7CYvEsG3Z2yl8bxovl499ntKSgy+95yTMTMnNyeI9/5E13Xn
DW+5XSzPrsJhgBy+Ie20e6MjTZeStoE8OiwkEmAVHJyNd8lsd/l6PSNOQKrI2kf2QBlDv8Mwx06w
2jgbSFbRuxE+SJXNkLxi4pile6TclkjcPlqawQZoEOMSR9OvVAeDuG1QsK1Wl2fbo7OebcKVCC+4
YOTR+LgbHdURvPd54EM9eg0jFbm+bmq8RbcPOZpZFoV/lMjLZcW4D2sjRhV6ts/OEb0ACeOenqXK
g4RdW3ZF5WnpRAQutA4+5p3KT83yfYf/VcW4HqvJW9nLkngAnnHhUtTB4osBaua/L2jf1rlUAf27
DrUwJ/f4nBi2V4H431TT4eUEmSJ43BP21reQzovaAZZXSKIsxD330ygJOLh1jV0PBWUBkjcEM94h
nnmvIu7u/pXafEpBSizON3SFJrzjgPy5qWrfcmo59iCa0sqG4nw22aU3xgaGX/U2cavKGATP4Qdz
v2qi155bKrgg7ZXeBu3w66Q4nmJIptcRB2m7T05X9LnkjhcJj07pyZGp0UPtKib16ZKUlia4vEjU
iYQBxhlSR4vWrZ/F/xFhp7VAR2Ri2VaA0K3Y9Y9/ndZS0aBjWxmKokNLWH7tZHHHjobCgR/zKGry
OgryW/Gh+ZEXnejc/7LSUHbQ5EBxSKV/xlWV2+lOPQVKC31fNWgIDhPRtF/ih3PEjjWxWgHJ42q3
sWs+x39INoc4aPV9+qBL3JzTN31bwMP9ckHhCuNiUAJMxR1Mjoy+emPsUCWx8to4pObEfCYLjVXD
MIH1FW15tTboOcszbzJeTSLnb+SVT7e6aEwuUIkpcZPsEsdKVisPDtg2FnKup2txFv6bNmkNx/MG
7EU4ze6K9dMLKh2UzZ1edDk7P2aORKGrbFuq9DO0rImJookvj3x06X66RgYb/u53O4HC1+66BkQp
JswaTo8XRSYN/INJ8s6UiPs1PmcvXWx0IqNAJR0htkdpKjUufVWM0hgcVj8ErdwqQqtulmhv8BcK
lEpEIYincWXjC22gEgrQe9mp89feZLdzHak+wDYUkT7DM2hPuJBR/3rlBYMGHwuPBSXPemL/jB3q
WovUn5tO5pc3OwN9G3YXuMzx2vDlukIKV/jBEGdSlHoleEO/5hoFBzm5Scqy0zphrlRNs3puZKoE
8Ve9HfjAX7F+a3KB4TAzkOf1Pbjfc+3WEXcv8f2bJzi5gMjpP75M3KXChuaL+lEAEtPRKUp90z0E
gpvwawvRZvA+uoqGg+j31I5UJ7zFT23rwKLxFKIFbb6iWoFxgjsfN+PZroXytjCOeflsPtmxjsV7
qXMFuvy1WGkfaBLH2sGmDch2JomY42Eka70zan8DRYCbUSu55lsWJRTWlg+VlLRoxHivVC1XDmfe
k5sZsO/ouJ+5gS1yuvC3rKeToTTfUaaYsFXgI1AyfWpkpGtt02nBg+PYQ3ERS8Te6xQhi0dazElq
CdlWkvuHGJ7ePHsvBpUKVjC0VnUuXeslIUxkaJbFO7terhn4G+xRHyL5xN2nQsoLXpCLiEIn6fv2
AGKUccCZkrHr7RaRg4Lj4XFxYrBouJPYHsal+OKp2M6pZlv+aBOrLA/qyNntIbu76qgMR2WNkJYH
ysyEW5vc9bbX19kZbwYDrWDTGhpg+iRN5rcbUV+LtUcHsfB5bj20uZ9h/EwJrUHH0kyAr0vpC1hK
5rm0gocnzYv0znK5XrS0dhZRnTKYDuzNoqgOVxQcLptNqHIg1HKS5KVIq4Q+VYT1JwFSBl7O8sh4
HcixrmH/zwBkNpQvlu831JmPRGLmw9R7Ok+N2IOOowrfOK7ygUesobVSPN/qKPNclHc4t4FeFoSN
YefVKFbdcLbshcGcN6HQgfcEkZjzM9ss1z2BP+szkJp1GYUemakCH6Gm6cxOhA0J/R/+lGeMqXj/
momXFwpCHcAqtCd3bun6yCtXZo20uSTZjDCwKYs3H4V6cUSGSbZgwKxGE00xGHizrzqU1lzhGNDg
8Jq0C6bZ+IiLieroKdTUBoXYOSAwavGieeIJ3yFeTp8FWqJokaqq2/hmnWh/l/B023czIW4LOxyK
LpnV1QxTnnIw8On3WtONU+3Xc3O+asGpEeL1H6eaGQxn+mXt9Qk8SN0zkmhSU8PIZFt0VYyKy8mo
jfYk1dOejh0hIBoPNz9i+cLFqz5krlV+Y6oIieMFVcwUujtjOphitIS8LyCdtKAvgisPQ+gYQfh0
mU7U72wHa4cKDcbNu2rcmOgvi7kMuc5K3VegSwix/a6uDJru2CvXkkHPLq3ZugD25DTJdgrPsoba
XUINlECb9YRDYc9YPT8+Wns+OZ7C7GUFwy3aqBGWP9jDThfR9p0H+7RCA+KmYeYnNX176JFrBubi
95Ys8jI8ijiGsHBKEIyDwZfDrfM2La4Y8bUNiuxQEny+LEj9/28blyO/JiLbGywp6avBXElEue+F
VNQd3VosCO5SbcCZeIABS7jH9o7zdlfN+8qwrCjalMZPhZw/9tEzRLlzdoJyDfUd164HRQQv0aoJ
qeRCsXnovP3fTmuOWH1v0M5NtCFjiwP71BvCKc2+xBhkFyn6nPKgFF5fpUXvFu1JA4kcS5aE2Zfa
HQf0/kC8uZxDOXNlwp0p8rkhSCOamnvMaf4Sow8O+2iJ0QrS/M7a7tI9kDLfk8sjb+H8Diayh8HW
vgtiQG9v+OGC3r5gvRnsjKUm5SxzwAGf4x4LVpM54IfcJaN16SKf1fdhY1ohcfXk5kTDpBv9gE73
yljvX17lAc4587EKwVNWw1YRG8VxDLaH+dSef7x67SP+D/MFC0IxYdcLdumSvoZRhnHjwr6RZUe0
PCFQcAg1eX+8PxYR2ylNdJ4w1q+fB/inG6qAxqFNQkBbcB+AdEjUEECz31GkBBuUpuYBs3NDzrC3
/qn8xqsCJTDVgIKXQBY0+uBylNI3X2rTKU1WQiV7bmcDuXvVI2Mz34dDkb1syN/O3j2TDlD47THd
Cw7WzHVCvpsCu9RjIA6xuXaZjCG+mlwXNbz1NPiHYVfCCbhnAgD3WT6wrRi/wavTfHYm4mRMh0Fn
fr/30EJsVddDLw5dyN0eHDmoDXKhcBCCnfkg52bLefu9X709jolG0g4EkYOyfRydJyMPTnbwfk6J
vzhiY5u0Da2gxMR/ndxT2kvLRdQ5F4RJY3nwxjTGVWl+cnYiBIkGnf1nasEI6AS6i7N+cpETmfH/
ceI3s2YRhJJFarslPJC2aNO8Zlynuq6l8Quu3i7tsZmyL0s2HeFANiADirNeK7zl3s8W0eVRJNVe
N6CTI73Ar1KnS60Xd/FBHNfK5XOruBV0oqfDQhEzbT1NQxDx8fFfgEwe5jnLAsMrCVZXxqbpZ+1C
DsMrXdmnHNpLJR//7y+45+9NXOGFGAz83nojmQaj/G4ilGLIUmMsxKji+WZ8qbWI/Qyey/IN/hYl
umSbaHMiG9wFg8FOXFOeQlp/gx+UTi1bGU9jog5M+dM7liJlQnsWrynbwORBK5BYq5IAbPrnmJ91
9L/+C+EBLTDj6koC3egRL4bYXuDgK5JX7KOXiexjx/AJ6Ss//L55H01Hri9kri668z4FFa7JhFml
ktKYI527jU4p1lCsE2oXmZzq2jRAZ0wsgHJBGackqkscEnRcO4n+YRRua8JpN2x9TtF0C0srPeyu
14PeZqmWJPHJUp9A74soa10tNWOFQw50zbX2a4plCKT6KQOwkb9dhnKovpKSpbojmsq3tVP7J6Vj
9qj3Vh/0eK4i2w6oZJRnMERWJHTy7F+mmzJqjiJQFqatWE4dCEygKie5W8SuNWYbmrgQUDPP4BrC
cAU9h9gLztj/KrV4PhvZtHNmpiiCVgCQdUNpD0jNrYM59laTFLs+4T5Mq4oyCwe0o2JiHqndPNEp
05HdpeewJcpNQ9ZLYBlfOkBXV+P2IvTqqpbqY9TyxZ8DwsTWkvHvi1qWMH3bPBKSzF2KnK7YlSVQ
Krlj1DUZcl4GhAn26SX4g/QKPytafIENOZAQ6puAsfyKSsGR8X3lfz3JuLDn+SdmKMFH5xx4xgv8
trmC3bBfaOdJa9VW7BxCuayTkn6sQzhQzOXODQMNNMvHSqzNGI9xEJy8uNgKuebl4nNrQwRvDV6L
VBd9Yo6IyvJtDJCCJ8XuB9muRQCP3ZNSe5FJpg/QID6VJmPpR74LUYXwvJuUOSaU8lu2YEsTUZYa
AFESxGgMZ8p56lo+E/yDffcWD0GbDD06DPlrGzYj8uwmqhmaGzzgJRU3/aOv0Nm3HaT9/tCXixdG
bFnZNEyRtrBJ6P4n0P6wiAxpJ1rM6iyAypY5NpN1wL7tsx1eGHWKrzN3vZJ/sRW1wiY6VmWQdLx9
l6ypAUwk/8kKH6UJxtWRg9ehOh022e0O8q0SV+/NaJN6Hg8TpzVVpDR0dRP15QhoVuKafPEk9hBW
1afgEx70XV7G+O5hENR5QR1JPHt3hK8IziVqKDXqhRETy8WiMrODiwexQX8+MdmsxTdXzIIEEhZx
6A5iTglFFTGOOzoYE6XTo6FtFtdoGIwSWlS6n6UcdvyR++85BwOuj6S3Z4XXLdfVfs+0NDMUnBIG
PQlNOrg3U/BgTnrmGEzcK0KQyUek0qkfapkK8l7mEQEbhd6Ii0Yj9oFK1Sdp4VnfCS9GL8YuQadG
s5yHxT7PjGjhhQA4LjexSPf/BIipMLNssgzCl9o7/zrZOjW5xNVaeQx9Z3vLw34QsG4NkptMGabp
NRj8EN/6EbPQIuVOrn+DoMuCw6+Vs6pTyjqt46rR2SI1jt3EFlnI5gWEEHsbrjhrxLtV2p4GyPWe
0TO5HinIqFl+jOcykw6hkR/UQ1O+Suu34caBrwEVmF1L9fP+fX3VzrdUTghbSTI7Lcxc1yAfyMSK
8ufgW2Ne0fGOjvD6cwTt9HBCqGPzm1zbHmWivT89hln9Rn93oP8EQ4sR1PSybbJl4bTCaelYXpT+
IsjffriSJgUCeoSRIpPsS2565GKCd+i5jNAV6g0ROPu3B6IA98v1KSqMRwxJ1+DPx1dPdrwZ8H9o
7iCUlmlI+ckFbzCWQiBV6P6+/mlGedxOeH0T65JDpC6ol2baynz0Bg6UbgHnItsNmsOrg/9wThJ5
YJH0XFC7XRv4o8s4/c9y8fa5zqQHRJ/i0lp6O5tKNuvdOGd9vC9UBN22srOQqUCWVLL8ob7T0rv8
wEWaIW29f2Y9ohTXSm97FW71ov3Dyfvnfoz4QNT4/v5byFLI06PAg4hdvtijFcwAzgYRtOlE57Nr
moXqq7AodnP4387ZQuRW/5eXrQCjcRC798RatbF0FbwtflPgd1tVoxiY+cKpqMv5AV0FDpzJ68mH
3hAd3sBHErgJV/BpgM5IqQifYvkfIjO34ZoL+7q24NtYhC+uthBsSF8tDVy2DBKRmPI+AEx4H90f
kHO4IMe86Gdq7jxAn5j5CMAn8rov/QeViO0PqDnNP6sF+fbtvQOimzo98scwIJX8beryXokRQAGj
PSUax0rXelRwxXq3r9iMmnBYV2es3q10/rsMpQ6XSTv/0q428x+qRTm1b1cIjJYYLaMMzGqrMSmI
BqZnCbD4scEvPF0+aRje4bzlUCwEo0r562DvfYjO2BEMovWGaygkxeUiNssbiy6rmBi7DLPvtJgf
fX7f/VCq5E+h7DUxHDM38pRlxFtzYbKGxVJDseo6xrRUofyB7CuJsLHfnnAXAPWp5XQaLihgsJdm
pQvkCe9TfhlxaxQEhEnaNXrtvSzgHFzSoSVLsnMCrUGKmzAatPftXGffSojoSdDVqi5P2KLkg1op
j1fXiWnMqFIowM7TRNAeV8Z3VdMhZ2H1LAqIEtT+wKX4XkTqjMulz3naKwJRk41MlN1wSRmTxwPx
J2zoqKnNs70p7Oho5mOEtw+i6WkfENqG0nVf5kNXWglr3xdIVVexp2CgeCohympBJVfwQBTPFY5c
mEcJ/+J3OSKQnRXAlWHlPc5RiB6WXeyqWV9Mp/IiqmQRIzSV1WQhni9Ix0dUpEpeW5RJHax5eS/p
PUjzmyLLfi0ZPtyMy3dXgpsFguyF8pLzE+usdR/aHF6MywJ5d5dc9mVKrob9mKg7fSjbvc8oeLRZ
MXC3V3RWw72osZvANOPo7BvlhwPMVONSVs9ARoAgRslIKdzJmRBjNyaDrSipnY9te33spvbLZ9tg
pq2k4LSFQ8X6mLGMI1KoAVzC/UfofOGkCmrZj/pbc1Dyvf0THL3mE9AEgmSZXsJo9p5U2svfaJGE
cveZzwf5WSzYMqmADk9kasfEC31djBZfaVxT0E/wuO+t2XIgcHuuJau/TfNCT749jFxu03Rgtpj9
F2E6Y5jT/+rZFx9O9Qg9Yz7Xcz9NtrS0m3BjDRzftCpx0QrSFqVEikz3m+vbbD6oZlqBnK+M3eZ0
V+OTh3gdgLFX61PlSYtYn6y/UVa0FictYhcS2m/LZPHem1lFrp+UnsE8odzsOoLxXT0bD/cpAnxE
sOGMQQyTYDTmNILsVo81f9m1kkjSnfNPszls6neaP2UdcK/4p865ddYJN2TINbX0vguDVmfbqBip
o6rk217P396yDZ2zWSVujupO1W49cKQz7WEJx/G/ADlHeysuFfYv8E6DlaSQV8B15fS4ApjdHA4l
5ZM+QISxlv45aHSDDLa/QGnGNYA5bR9tA3QHzEWyrF3w8oA+w8U4+7LQLF5OzYdmdWhhckFBeGrx
/FEYAe8PKh41ZU1PvIOQ9fTgQrgrpctvkLk+Y4xnqXFLB27Zbp/CAIPWE2x93NiQ7CVLAtxiQIq5
FR/MN49YeUSimXHoY9koIzhRZE0VJRTrngfHMvfvFsxRwtvY0DqhjVoXFzqtwt0rYdaXNVCAJUkF
amVV2njbOLAmElH4uX/mVUqpT44qn3uSRJzlmlsZrXQM8g2gb2v9wU/h7eGfUAfEt2J7a2lVtA/X
zobSgd+chj8V64mCzM0sv7XME6rbPeOpPyz8rgcdUa20lRIdUHKldqpLudtH4DXIO9B+RJvpAPZ0
PHUzJIAOBkaEcSYQ6A6ihLVzm8eJSkK695zV+7o9icyFjYvpG3z3T0MlHiBRGK2hOjejF2274LIk
vVItULl41EANSIaiafsnXN+CHN/SXyfjWt4XwIPZNazeS8UBauHzWtfMOliIDw7dAvrB4ZRZRJ4n
kqLUwdH/cNKAbS25YSoHSur5B4JhNY2GXuQNx4slbpKy0A8Wpdk61eVHEe+wvvm7poEyWw/q2hde
nexhhUqFheCA17Oo5MjeqTzAFzgcZzBRevQsILXPGv5UJ3RVYaNHALH5AboEBZdva21uS7P1Zf9r
VBvHEnT0qPjazlKXcrcKiz/inrrO7FO9if9JWVY3lR4mDXRdNXHXO1/ztuQoKhtjruWKvHGQwimZ
xPEq+SsGPQjxvxguiZb6+ikk2MYW5FNjUONArZ1lU+WhZtS+nd+GoPhNuoPoIQiX9jWEdPwWeVca
dN9NEMaVxmtrOBnD0A6NahowElljR/Vm6Lq71djjf1r1ETBNiw1BxQkpIhTEqzI0JiJa5yu21R6K
8S7DYPeuyiR4vVkbmWi3U9Wr/u5jfGZB6dv5eA9YtXa/s9cM4UNQ3ZsKmxOzPVCfpcSHl/1jcvI+
lLCRqfvXCJdyCB1LSZyYfXXOLY67R+3iWRFlyJQjo101I7Pj3v7bnooKH+46h8tZ/AYOFEhoUJOZ
GJA8O3rk1oxwKZDngUTy6V+3FZsSuqsjD8UiCztaKV/KNxjO2ikmkMRlktpEe48nRS+X5ny88kEu
882RhNf2cYdZc/Y5IKtdCQw4Oo8529N00rXPFI90gCqbRu4Lf2uAAvd4zzz/8PH8saBCYRjm1+h3
N7Jr9Uqohn4OTze+6c31pkGq043A5V2B4Ww1q77WWA68Uj0ZeWLs0SKtJvH4O8Wp91hlrEchXz5H
HsBprg0R+jpAkX8itSH+ZuULNWM7eHrOArXczxT8kPmbCx7rYSRpK0EI9Pxmk9IaXRmNlxvnzq7F
zw+WQuIF1RnFOaDkFn959y8dOV6rifz3egltwhBt/m7dg7zf9vhhOiqqhHeS2/tALMXjUSeSwHTE
mhgzjtGzIX7xTv/bJvidpEimSN9Yn7zEzVv7uFiGGx4veZH0ESFq0fAz3UlaW7UfOzkHDOe2qGRL
uxmS73l+IMEzSJ/pk7biDyLBXVCmy75IuI8Kw1fJ9mE9PNLy/ZAV/GV0yLrV3EAol1aL3hNfWM4P
/AYey3tnq8/vq83LwDCkU+TzKCCUXxqh6/RkyZmZzWnKVp2j+R3HHRubi8aSaQkcXENSL5sxE8ll
xXQGeMktXm6/AfsW3MKBmn1ECS+hHyHSYUGRLPT3214JIs0kWca4pZc+VTQKw+QKlFgQZZEQ60og
gnjHov6E0PooZGNaJP6H6bRu96AQ2wIRGhlJsHRVKC/9WjDs1Ax7lcqze0aGrT1vyNt0SVCpE9M9
9ou1x4e8cKdzRSyyOHQi9lpswL25+S8GheoVLs7YEP9DK4XjPsY5ZDBeebeMXlv9Yon8uKgrSDwk
u6ZYfodrEDU4IlCzPu6XC3Gy101ZsGnt6M4x96RmEBIGap6alhAA9ePlLFNo+YiTkcp2qVCOSP4i
/PyI+9/oOZGVnLtGh66kzAsTLskQM1tL+ylGl//vRrv8PSIt374Kz++aZ3nKIYx4jVQ1NIOwb5rL
w9Br4QSB8ZPlGhC2L4lL5QV/AQCeOzk7kVUunistj4XbMmSrabiGrGW8UOX5Ks80BjeCu7KYqrh1
u/pphT+BKfT4mCUP1MexRRL2Z52JDG9zqQdxhT8TLbNYAfyR2WOpCw+vbWw26swzpNJ6T0zYFPJc
jOKTPHyMe0Bu6IGcr9u3DwqYwM26pBwHH49YTsVNm/N2DFqH57dj6AwEnBE3xLTFXSF2xq8nOgC0
F5uiP03JQbJCiNFhJz7jfMOzvXWecvQ3zFPN8oSHpxs/ODR9t7KHaNXZeBA7x2oPExw8Rt+/Zxtl
BOXCWHiPNEkgYDJztsgK43HQbigaRsnrLtr/OVjuWR1MoH5ra9F8yc64WEJ5fIqesYr7/nLp2ywY
aH2ukMnKke79esypxD+afmAETIWGVoPgGXVsxHALzmJcd4X7Pb0hqiSFBpKG1fvnz8hGDS1WlwMo
i/OYRuVGTm/rV12it0Z4giexuHTt9wASdYWMzsWmNqzvnmD5wh8Xce+elwqPaDXpcmvWtzcrlcl2
QlqfPCu11AFQMqmNA//eLVx4cZbuD1BmtYHHIJjwEr4FDYD+hPfe7T2xoZsZGYp/iRvVS47mB5e1
MdYVEfM+ASehJdKl0OcM6J8yX0CGW2bzL9MeoehQbDoUMJGmveNQBERy5KWz2PvZN3ZK6kgYNyWY
LqAARyZWrSXnS/jtPP4ZsaGZ94WWXliEjSdVJcRaAxpQg3gnnVed3nBN3oKsa/CFirfSC08XppTv
mKgVZ2E/Vj1m+UPfpnzw64JJGi+z2a8aJSEbrbEzWCLq67cE/Zpi2UM0eNTzZHADzp23i8rKgkVv
GbIUNhK50VdWPGgz7PHDf4sQc79W6eo2Veq8upievKNOrMrDvTCT71lJ8cBIt3ZlnDTl9ur3WmF4
fg8j48fjIOfQNGKC1vIIPG8weWXz2n44VNoDHDlPNv5CMf6vrRBxuImIshlJilZYyiAHkNvcVCaT
m4Lxrt1O0HF4tGQ1Msa5pp7zddOTG1mqiWyvQMqWZHhJpE4lfHVXh8iVRGpTHFs0d2RE+WQGT1En
GZEPu1gHgQ1+bZlF+zgafDOd7PNRzoHv3xr3CpjgoQD0ybRmjcyXxWTjwqAs0YScqauf2ML4kHCf
RTiznaJPZdr6tw0Dh0r72GRm5akv6UvXQPquqxeBnZJFConJUQvqi0PgIaFvnM/fIsA81qN1nyUE
5Uz9TiEu0vHAf8EL5Equw1MjfdXLpHQvuHI/F7fgSDwwTv4bc9oF/Kfo4qGQGM/96Dkz0EJOsPH9
i5+a7BgigQjnH/SNx0RN+F3R6opegTBos0B+lDzaJkQEnF8aK37RDaeSee3PSn3Aj4TmKZWoYDCR
M1a3XOrPkTyEgtAByHKkeujuOKEo4T/NDh1MpKzjB9BTTW7L7bG7HO4C9Usl7+d1wcy7XyeFwhiD
EtaZsDzvlOU9w315xILrEKY1jEzapBk1blxd9tCTZxJidPSLfHd0FgEZuNRocrmrBxiw6IHfAxkR
wMSiSiqQU3gCG7Vt9hv1tfiTIPThQnfPywCi0ePNCGKxmyxWht/KYfhLm1i9rJlr/0xRYoD1zY6B
cKjRHJ5Qaem31n3sVnICBBtjifLqnhWJ5+anQ2n5lY5YPbdFDw8HWBp2fjL4rxi7Z8+mOYtJP1Td
qLW/f6xE5XI3pHez8pyIE+J2vN41SmeP56o2yLUIXDPXtahVgNvVokWO9FykEP7IvnCO9lRTmhfY
Vtk51VUrbI1nSXyg0oIcsTe9CqNsAKp4VVxwpwr1F6CvjeUJotFZEmA3O6P4eY4AJhAzMLv0HY9f
kDmzKJP/1l8kQj1tdMrkAX/c6rLP0AUFLuzKpIuK2fNpLx8hlEp79y/IZ2jUMGYpvVv1DWKSKbVo
8/g+cGKgl3p9Rkhm3qrAkTdoKEDuF6VOcmq6zvQbkNyVmiSDVsIc/jEVqx5NAzES6kldxySftYZm
g/BtnfLS22PdADngrHgkvvnQj1/nMGZM5BHCH0mfo+KoIvmC70281u+PTcXQCrYAJyAixcqK8fLN
fndcnaiwgWIHId0G5j9e+u0L8+CpFcXfwE4FM8AIGrrOMgueUQ4UOyQqierwLpcvlZcN8gJeLXd+
HX/0CFYtr20zVh3XAtA94IQemH/3BdkNRmloUOp6HWJopd+AffdnMnQNZUpQNGKonrpnLnPD77uA
d6JqQYa6CdJNPzXlHxbalW+uxyNniawZsiHCMr/p1WzttsHkLFvzFgRJt/LzVb1dTzEKoUheLEj+
x9khLA82bG+/uO1Htpg3zRuE39tEDHF0d/cjya8BYR4swJwBlqSbU7vUCMCm+8hqnEXOiYoc/e72
ymso8R4JliqWAYxGk40a2ng8nUocmI3SNCKT2dM=
`protect end_protected
