`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
f/HeBIsD2CdoDuL9Ccw4w6DLuPNmcnZIDePd31zo/fv/5szwPwrYz3j+XlJ0PMRkgX4zKnZZ9BDa
h5Y2tj6HYg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aWIq6V7Jb8q9AC6TuGLPe33l4Y8OGFr7Ar+4JkdgcO51jetE/cKNkT2dOcPnIN+unBNs7bQOKf2F
KqaqLXTzduJ12hwNAV50Grvjo+xTQougnOk6nxrHrfa37Dert+SKsUX0b8hNXBpTdDJYU05gbnv1
aLzZcrRX0boRp4Mo6V8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cedKQpTrLYbiYZcy0RuT3jzbmuz9I7qQmmpAFdzbj/eJlguOPHiGgSiH+54VxpYK55SFjtvvs+Zb
WUgQe4Vhz9Lsp/j4JuP42MVWwcmwetlxw7Jp4MUvLTuAnTejlQKrHKD5AjnAihfGKRDTToAbO5HH
pdYx2nBrWK6CF399ZccXDuMBqPI3gRnaDaLEyb53uCmlZsSB864zm1ma2DB263r3CA9GDPQNN20Z
7AA0aK6r46kpdfaoGdV9xKiQtGYerFvZFw/UAVNkzh7wJi844mINuLAVMdkKEyRJ335RJlTOrmGZ
RE9Zh8cLrdSqztBWnV4mu1Dn8uJgySSnOXRePw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PsTx0i6PWL6lnB2sx8EAAVS74eThqWV+/zRyID8XXjR3gPWs1QLHzB4sqEv/jrIJI2RDBclzz/ew
mKK7EGxA1az27NJDTzmGU35OLDZ3SgdNmMZqobKEXu/l7CEo78kga9BESYaJEEOW+vcf0VnSZ1ZA
7ubZ+PX0DlfnZCnKkeY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
00tG2Ar0TeNo8dxARfREqI56ra3FCaw6SyHOrONQMBCm4YOPj8STYCPCRQUAhav9zKE/sTWa18nF
sGdejBdSDxOwWM4xZfj7YGjOtzMm/G+7n8SNwrdCnFJKi7MEiodUGta1nqmCeH47/u7h/C610lgL
gxj86R4v6d2Q8yu1cHvIXa9GmTs2fZVsdNJ6ICpe9y5/7KykZ2X17/s+FYXdEY+g+s7fNkW/5NC9
6lYEyL6BZ6ltqzP6L6FZCFHj6/R75rfaY9ntt+CIcqVGW+tGnj3+JAF2F/DNm/NXj3uLw6J0LkR4
OWvwsDb6/R/QDIZYxVCC7DHahg6q/v8iwSmZeg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BaCQ+xbQ1kuC+RCKxxJhXlSfCvarc4dkeXveWmiiPMq3mpLrM8vRDX8siy05G4jp4tMcup9SA1FD
rOLiHIWsVvK4NITV2dA95S6Q7PDa3n1Su2umzgc2v4tJVCjM4PifdhWWyEmzjechFzf1jxQNe/TG
WQpSbxRjQqej1UoSj4YKLgvJKBeKQJKW56i4iDj2I1L9Nun9elyVjEeNdXAcsevJlRdaorB3vmzp
89beYHgk1H9ftCvFzcgkl/jF68VxKnAcodOi9/Yo27j0LwIo+71YqC53ujzpA+GMIoCO0g0/3aYT
KHf043su0VfxgNaBZJvFipTcZ6o3fDtfPgAOHg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12640)
`protect data_block
ccZm5b9fXQtRCnuHWixUNkTAaXSsDd6iLm82DwipjImJnwqZodSI2w6Yxnkg1Khg+OpsnDNI6TAw
ut3E6+AJF54jKzYJf8Jc+rUF/62dm2yXcCei5J2kHqRyCQIULuWpCcpBq41GhUXUZbobyChh+mmY
RtE+nGFyePW0C1qOUNOrt8A1cf9CQSU0L9laB4f0Xv8bw0KmTrtvl0Br563mPURr/4etowlwK71v
C9PkEN6ud6oGHwW+V4mFQOnp2vMn2k/ysmiBH40PPWPVNq0n+qvcz8026gW1CxVmGW4og+nKHus2
e3BVmiutL7sdXDR+kO5sBt1TV3Ga8gg5TzH1J32brInbKtrNMgqoZGA47ZZUS+v1uH6LXH9qXO0S
ruVqBUJSFxhHLfAaqJWPVBzpCv7IvMoPmeT8UA4+YjFWyyaX5SPvyqjB705SrNJxDz6dtb53Qa2/
3hPJJZmRTBp3ocbneklN1D2i6p0azMtT1CWe1Lao8+Sp8fWmLoTc2xvR31/Lk2auIeMwG9kJfIOa
rODU6gx3IDf7bJ+TFTt669YxVKwt/Ipmrg/R0s6cyxizmaPoHm9tgwGWEoqUIrl89ZSb5/UlFoyZ
qedbD9eUjr+rRY+ly+fBSLJR7ZqbaF1lI5XfyfUlNcFAaj7Gvvvor3aNVvHyqtjExxsmY42V5sg5
NZFN7psFLdmVnSZfje7xVLWVnoRnXJAUPX9y5H0RhOydSj56QIhA3GSmcLW4gDdVcwsKBhWLwLEr
vxdqP8cMVHq7xVoioJtbqnm1V+qFKmVTXLA0sOHS1H22lmJuu8A2nL6jsGjJao8kZNsxoXEUI0on
TODRrFur5H5kHKyZjZY/kkDXmvU7yYsWdao3GHQD0Un1ghH1+lFKps+pmg+qSFcVD5EI4guTLo7N
3xC97bLDtlETDe2V8SOUYLPLDnfCp2O634iJqSs13xVfmMs/3b3VhzRI3hmYPMrEmeCcovjvfn6C
hJwhBGFjPGLc2Pobz158dFwyTrTuqoyrfRdZl3x4pr98ZcK1tZ0gQ4RA3YI5+yQbBkKPKEsRiEis
sjbmUw8W06uS8CTtFZRCecR4GCtNoLaTKo8AKyzCXtDq6NLzN2hbAKJp7E1WZs/kV+6G7uICwmq/
s71eur3OymIzf9rYvTFx+ALETRQi+zaWtNxh2wRFocF9Gaxd1F+fKbujj7y5PfN1fh/bwMY7Z84C
Z1UmdMwd0BchBEPhcChyICndnb30hh1xarAbF4p3MIug5/G/ZUDb/CitaqcDmY68NxjWdWdP3f/9
WcTpa3o0dCm0V8wTsjr92+n0qfsDrSHc7IXK7vY2qQCF9e2VNm92vpYAo9FQPLxTaIv04ZpX3kHP
PllGNRLV80ajdfjSmXp24oIA2s9vz76IK6wNeTv0e7jGrXijF7ag5P8cxrbj3cqe6BdWl/9jj3eT
7Uww7YVmIcS0Qzxy+o4qH9XqW/rPKgRo8bQpFNWxU8VEMGanQw0ulU/jK5fQdKN1tnZ14dXv6Akt
SaoBnKJFWUY9B7fcrBeS+F8cRmU9wJmzQc/hngabOjJdmV352ebXzHa3XHAOuEWkVMq2Ljxzn6kZ
8nfrXXW8qwdkgGbS4u9+mBL0kJLdGNLpLCUhScWvRjujzsQrVuxbgSePkp0D+6jx8OlUhN7Dn0Wa
od8EbGHHDjJo7XJtGW6Pq/vrdFRRFy0Nm3UHwjyfuNGNzERiey5omzqVXUXX2Twd5VDD7Ofgjzvl
Y2XOo4BPlf/5EuSJsmZu6E8gGTZIRGztFi5GgGPIYwreL/IRV7G2msKTXpmhwmmNl8+L+Q6uhzP1
y4OB3MhwOfbRuIEROxfydC8kz7LsJ+04Qx08cCTRccCEUGW3rLxC/kTUN/SqtPk/gRfl9A0mEvgQ
phuo+gLfTTrCprQM899dvveP3I14zwYLIA8eR8OfacsZjzS1+lycja+6P+QyFPg5GnUgxg4p9E1n
fvWT0hdXPiV7rTqlPau6/VGpGYynEPbEKhxUc/xvAh66vYQDjUw0AFtRfkqQoc+rzDSn48YVGBhv
zQlgtrqx6qB2GdGnOdCl4C3ZMyCVW1Pm8P9oI6GOBjbTCOoIjxIpzO39LXIiOMzdmEdXESYgZyB/
fzPUy9eQoCK65TQ+KcrV1NQgIx4+hlv0Beyu2RdGkz0Z1NcJPEzrLPah4qaKVQLBJfbRNqOgFFxB
z3cWKOz0SkGDuaz+yZT8a2QslWfdDRYQxpt34fy3TcHtlKu0gmfKEt5Io3YjWCV6JoecTUshuQpI
33351Sx+YNch4D+BVOY6jR6u59UtMm/jHICPHf44XdPY8UYt3GWHX5Y+UQYvlMxd9cmU0Xi4InEn
D0H7FWCb0qA3IiO1Z26ho1oh8vcGweqPBUH5qg4fxABuklqZuXZxwveYcM6s9KzudwHPg4KXHCXb
MuFRSdyjzlvitWTKvLvJK6niblVaIEqV8eI7oEx2ot6wCCgdjxhccHo9UQmoq/2P2cbZQjxBiXJb
5jSYa0eRXMsBTQ+ZSBQJIlF6L+HrJ1md5QnNJ0jgVsjQoWHAzcD7G4ti+k6NvETzr1Bqn7u3ciES
Kd0uNSkfEUE7h73EwamKAV3O0P5vWYCn43Dd37re0EfRJiuUdScQneGwjus1bgK9kCtIflbX/Tr2
uE7zg0OpgLLucJPQ3SLEB7LQbwx23HJRHryv30MUfwgHBuxQ1UfNkpIsfT9rCXb37D/vDF/igDIt
O8kNDlJhru8bhKj6xeoN2NrCQGpEOKXWBbg+w5jkXAt9mGHx9mq34kCcnbW8MqYROFsmCV+nrRXi
3t7Z6J1Db38ndw3oqt/ERbeGV/bVSp5SF6tLxjfy686H5jyeTtaiftfQj566yhOA2PuyQSRHfnN1
mSoeFX6jWHMnPrr5PH+wa6SnD3hDkMZyc3JXM1Z/s/pBgsmxnLpY2SThBDPvGnap7nb4G8B0eQLw
xus5c1fAXWXG3qctVVWpvBKQXVSs3ieKXaXn8oCQRRLP6RINYsW91oFWmm/klRowM0ZJi7fVgfbe
7j7uI2IfL/C4Zjb6L/UiBHLRST0emVdr90UQ9GeMoifSIqeGqldv2Ohl7jgXJe2fDerWBJgOE3mi
4yxe+/eYOc4w1LW8CvTnFFYkDCboGMZtTfVFryQPHLztJ0mxAGbPBf89gHiP63ykf2PWwn3F0NPW
SkMJoxmgGF1Xzgd45AMBFGZ1DJaZat2Ljs0e1oK1s+0Lx/OQT6U7+pZqiZs9r11A0i2um9hvJeZL
uqMoz7kaInSYJfVuU6beXcOsq4PdwJ3uvKFm6j63RkNSMIuB31TsbrxqoCbT7KaMwBxNcTFSWos3
lBB0LKf47pufm7EQENX1OzSSgGcqespYQ85ehYfZ0krGAdD1d3S1wC5zkV0Nc9oPWRlNYHbvqQJw
X/6Pd0w5DLhYBxaUjOhjE4/fs1vJ2tJqrxtxP3DYEK0/LmbHX4aXgNjzzIgnxKdXdcSwfXO9Qwnt
RJeRU92id7OzggGtZQxMKMNRnwl2LZZGR5XSjqvBIcIESbUU/zNhYxqT3DvAEvrRF84w+L9NfBLi
hEi7YfT3TzzW3u6V5xwGorfiFXqygGj0ibDnJBqGldfzJhSVZRVSJ3/3NnCGLyo24p/Hl2YjPQ5i
lXl9TIwL7NBLvOMJa8aiiltfjw95ddi9uDbKGchFggrSsxxEd+15IjsC1ZScHpQs2snevztP5acL
G6YzDSrshvBWHUs+TP2AMLH5W97qinf0HBcjkgqCa9snwW9hDhb6NWc7R6qsMoYu/0s6BIfahdcF
4k4T8PCO6/vDe75wbYTbPfRWlzVAbfzpj+Kk2VYyM5Qy0N9/l3YvAktYkBiI1Fc1olq0tjSrCnb7
XOIweBj/thauel9ufp8JfWtW86zUx+y9UwMtsxUnRGCBkKjX3+3KeQBpf5bCzkwhJRENujiqy5YB
YH0a4KKpLZfOs5XbB1s5Yd54Y3qI1TFXI0nd3BlcySDdZ2EkehC8IU7u3iDEiiMl9hQ1UZAG/MOn
/W5okj209c3NBDeq54mPE41TGUK1/xYO/J3CBdS803iOVO64lGCBfNNI+RTpHrv9Ci1+igTxrn5b
7gR8HulFgDewIGoccyyhUjkjSg+KlEn5sjWMM+k+AW5SaitKgx+R34t7FQlshM8brVCqQVsO5EfV
yylwUcE/QL9mAZE7tsU0gCwxdcpPyTT6+3ZdnbmYGTT4i60VMqDtls17yZmFeG6d9rrcxGgM5Set
VbrVhB+lPPAIhUgRHbHeYrobip7kMl83i+SRnsFU5m6sy6MWxPZ1GMoAST1+XFqIlHO/GjGsaZUW
zlv3eMNJpK/dkNcu25z5AOjM/FpLiMIPidvA5vIMbwfZSKFMB9qsWMWy1JuA6+3n8MRf+osz+P+2
dql3VtuWe7vRdLrlYaNCuwvvgPFrO0fv8lqCvDGDMM7tEPH86GD5pYuIOoojL3tSD8lD2Q9JG4wS
71DKhjWXCuU5c1B3cOTZyyC6cicbRCFZEcCh2mUtMxDmxlGpDYcqd+QvSvbe2GUXSrJKsovcfQze
a1YP4eRgrv2PQdFmL6aTjHy9PQ/wzMIg5WTcp2kTjLv9557YALYe8Fw7w4YnRHe68XTkH3T+/JsW
/5aieBNqB1PO3Ol2aGbMRyff/jcS/s/1ixxzKnoDTjuD2qRTqc+t/RA4/9HZ0sub3LpjwELPPQVi
7SDlQEjizdCOys2xcOhA2gQYgI6Gdem2Yc3YPIzQ+E9lYnR3ZslIPTIrei7lgTCm8Q6c4dr9puv4
h+zj5tg3FCfOyDlHjW4jgsmvMoem0egrp/6dlH49mNJuhC1pp6TPSgZCLPZVtKvMVphlqm2v2HC+
MKHRh7X5zaH9Lk/sbWk7eUzROISuLFS5ZuejILriDPqCbHGhG1XCrDidGRfMh9Ib+iK4nR3dhLFu
//gdViaAf37dyjf88sLSRQOZMIyLlO6yq2V0Gv70IN2q+JkStBeKYj5KW5qUySBGqjECKrMzFza4
wfabS8WDa1yhVXWFT+QEiVKO8PYAqLssFDwI6dMSgNs9nZsH/LKDcBMtXbMCSou2J7rtZY7DS1Ty
1/2/xt7xootFZsp13Jp+uaAHYPccFVuMvRJmYgVHdO12/gl4ioEJdEiKaV8Ef8+L9uVOyihb4fAI
1ikhKyGZhEXkjy+CQxVaFUwGTC6uouQoZl6nIi2fWwtPBj6oAL60wIrpkDRZGGm7rhAzF61IGVbZ
4cUK7eoMw/eZV8X7LUz8fx++/tURFzOwCIoXf2n9veCluJ2qgLQojua2h5fmlMrgn/5O/Fv595q2
tn6rL7BXfL/moaamSBIGR007TfzZW+dUr1PzDnMIbO8cY7agYEPXLrSlmwdBEPHSbi38iE/Jb/Ix
qPWXGqVo5bt38VupemSiU4tw7J/xFV+3T20v+nH1lJKFzMBBbYmJvqu2W93DXLB/CJIop+uBmHh8
SI6oI/wMxo55AqB6X9iGN9Kg0mR+eJ2dQcOV4IQATAWqMWlszKxECbl+46OJ190kh24NzhW/xfSX
R9srAmuGQwoYeOSI8SSbDbySZGA51dqzUlNdYP0U0gLRQGB4xkip25AxFt1wpwlsVCbwI/XVE+GU
jQQS/lH4g/FashOdoJvirUqCj2kdw6XbzWJQZJuko/8mlyBuR+Qmw5u06bGeq0vvWJ3BqADY3+BL
2euco6FNC23GiY5rJfq5TYcJ/E6EXFkWV902gYX9N2ULe5WMbGhyu7PeLb7eiPWo7a8oMuOVKPph
Lo+AThSKqWfc1YP0l4bGkCNSjVi0QynLJlrhrRPjAthuXB+ZYxEFj7BtlkP8+o4XbsB/x+UMXrMQ
ZIM8NAOiR3KrhGR00wEf6i94O1TzwG+RyZJoLsrisDQS/3RBtyeEQz+tgrhSyNcI0uJD55gu9Zqb
xfCIt7Ruoy20FARNp6X7rs5FXloT3Tc986oYwxizm354uMqzcBWu6FO9C3rAyQi07lLgep/ftmqT
MZ8NwTn4dkoeAI34IXmhvjraP3e9o/5+ohIQ4W4dw48LihU8e80zCFqWhLB8bLWqt5OrIUVXMKuQ
6/xcoBLr0mQWKX5VDrnTZR8AwUnSEcgk/1XDiA/g9DxxzcvFfgrSKcFgMmj9Meae3b19ySVsNlHx
Ercv95Cj355AQjiBTHz6uWvZTg+uHBXEP80sBo1EG0haR6SC1QXujvTJrvnLKi45lvDsiGjNPaL4
dAh1q2TOZYsckQV0oxqK1o0FYB2bfQe1IwBccVAiu/ePCOcqr6AePiQ2DztTZ/hXFK6dYQn9a8nE
BCUrvD4AZ4MeAaT5nJYxlYK3L2B9cxJp9+TxBad9a0qQ99bA3EXa8vzJ3pBxmHkwrfCUYbsYFxwH
0AR2TrYD25q+7v38NTRkuI+6rPrqKv89RK7sNKCmqLdonR+JZ5am36WeuqJtdatp+UQ/H8zhe9YZ
c/wXx2IYPhcBJV7CvCjz6dNGUBp5wLAhqD6wpHnA7/MmQ+MGAKSxXU3xN+cZxLZemjzzZ/1u/3tA
XJa9TGhCaOI0fGkdTWeR/SCK+ZJsQrFEJj3LXKg2RPte9MDArT/L7RgcJz4VQMymGDB9Yfz5CXAB
dfTrTtoW0ejb+pBUY3VbdK3fVIXg3ozIapPB2sfsMZFO3lueCp1ngcwuhZLgY81OTbnY3+cqh/tw
pPZVhDFRr/3tzWxSKRKUyFM1GHtGzfdmYR/QwfjsZ1ev+5W9odHH91ZKMZQht+6l2Yp8d/QAa3BT
iEpwZGHHjkqn5c3Kf8QDhNpoAsHzQ75DaqcDgzWgn8v3ds78qJ/lPHAtLqMFoUxNaJWs89VzJB7E
CBKxcT8BHhvsJ8s1uRzZgv2UAx0Dlmt8xhyN3CaC1ocv5RwU85WY4GePs3XB2C16Ee5tyryGIKO3
jnOm8FkAewBRDj7zgCJC2tMVM5Z21N/rqI3zBrTsKjGFTOkwZ45+eg/s/FlZsJWeKzN8cp8NBGOv
RPgUuVly++PH8eo/c909t9a+qtd8sVhCTBG1psDoJ+aaZtkE1K474ciAsfmevyBZmjD+NAHotFIO
t7/m449wd5XSINnip09jfmSCO70wdrjFQ/PdbHLvdVoq9ey3Erbu03+y8aexLDq5PT6ip5eeG/xN
OWK7uIckYOVEm3/HQq0CLZ18iG1jK9lwu8puYi+HPmeMNt+y3I9f2TfV4asyPCflxJMfnTUjdaAY
fNYHpHnhx2ya9Qa6GMGaCmZquxeQynXr+DXEWAPvX2YNJGMRLOs1eMUJAT2oMl+W1dKuFL7wMALu
o1TqsN3FeRUimkddgxMeWGuNe4CRxYHc1Tz+qKu5sJj4WCJmHSv+46Mi2N50NXEa8qeHF8UwJYI/
YpcOrJa/5yawKPBi+pQZwDGV3ZhntoLY3tQvIYqq4twxYwzoQj9nTAvk2LBIhJzN9hHjjrFb1f3h
Qeo1nSCsrdruOVLHTuclp/zHnmkrFJiqhckE7RnQZXuh+K04op879QR790Cf/lpelleGMyArEiOr
pE/WJjwq+G+zSIDvdfJiVD1lUetBQzeE6+dA32pufxRSeAJoMx9Ya0y8tH/tLlkmjoB3tcqBcp2d
oWT7epcgcXSXDNng01KWCKG2UjUY374/NL80luwgHAaVA5nrNEZk9/fZeTU8umsab4+ih1v5IG7A
zDhpOysxUL+Lly5Oljg0QXjf/mNKJ2u2s1ePMxgKKIqcyNJ3YC3jM15fT8U3QbaumRbvIVn5vV5I
61IGB1sJtHRSrW0gRCvwAIbvfSp8lgK4NYzQ6IhD0FzOsfZTyjINUATk5vmt7rGk2/DxKZHc75aR
eurkXWjPhMfQx1XB0ZQmHRvN4grycPzE0dC+E0Sz5poZWCCq28AjryfoIbXndF39tgwZpg8wkZwH
b2r873OIgvXcbQZTM7kcmWdkod6F8Sqepka5ilMgUcLy3NY14PYRlmQh5WOCv9TDhjl8t9Jx/te5
PxIKN9psos/TcZQBzF80vrLZXjI6lOIu6p9F+rSOSuQsVaioZeIrKrnFADOJuiSf550EQtZZisa4
EfkIHiH4k9vtTgnqc2I1eBsC7vvDgVfmgrhOahyHfyUiS9W0UoZ0SpKP+us+v6GKYx+Di3O5oUUL
PrYns4Mcy0PrbTZ1O5TFLOq/8+Ufoz/8XEiohvFW6SHYnSGCuIo5LB2xIzAMy+CSJj06J/ZTelVn
v8IXQwjQUiHK1ZpZfpdqxYAe7hcqejOg0cK2rkoaBoki7f4mZOK0pozCnphKQ1WxIoM7EhKImyYR
nqvsNaPGrn3wdhWrHQhEFnze4GJ2kdXq08znmfkywX7HUyHOOI3NKysy7uJX+HuS4MvRyleR0WFd
BPVKqeVFVU5bzP3EcNg9P+79k6UrbLHUSuS5n/8L0w+2zKMyjpKxlj59/zYszsHJT5NKB2t6aaEf
xe5HW+ugmTWIiIUGmGHVPCqZS8LbMu91mpCs1nqELxgL1zKgs0yZD1VXW5t5qHBlrtEIH7nyjiwB
EJFCcPnnqsYXoews6f+4frlQ3soRd0gp8a1QMQC3gVGhksKb7QDmCShCmdsmZiUBFZY5IwCEGTmf
vvK/E+jR0KWgNgxkqN/WVQbH8T3SYYkMW11GYFmgnGdFA9wx9R9IWjS1CMULQhWc1ZwA6AbSDcSX
omx1ntzda7lAtyRxuP2wfSnchmi6UATp3iVLuVgjkDv8E38mg1pi/vqrJnjmHf7Oxq9J4tttRz9i
HSb9QUnhgGAc0SH4M7aWRV8V1zh2dMqKSTPySYGgX4kyiT9+JtbnXUQC4YY8TM1LyM/3Yxp0uW5E
awu6jFBW8/aBaWu7JYrQPFspQgF+30J2Qkqw7reNFMrwiqZjyuydrPtznfJTUEZIXZuLZeTZjU14
a522v38N6gx0DpxKLKcm5FrReaTHZQ4OLsKOZre1o/L0ZId1isqvMIKeOMFH8WNXggwuyHafxDz2
MbPiaFnzXcII9xl1stc6qqQXn6/pChm2lWp+oVX8i4pgbhSPGLSoqPnjiQg3jy4gERtuF+ptV/Im
QwvuVfprQWwjDusedmDLLV75qjoRncbCVBmngkMykqSzFTGudCSDwUwbaJFktzOL3HccPSvT5EFr
D/rnC8Z4PQyxrjuOlnh/vZKlTUBdtGS5QN53uPW/GM4hrddY6i1AZdRz/Kg0nEHZ7CqyGZelCRm2
kX1o7a2I55v6K7mX6h3ZfKgGdA19qCzLYC1wuMtSi/rgg5AILTNXXxTVggB6B9bpEcptLTX8/ITC
0CWvG4xlRt2+vxVqj5O97+cSOqAyM5cqJU+vOxxoFt4NGKVNNazeacpBaouJtFqFUtoH5esyuQ+2
c3U7sDjB/onWA9Ni8/ICYw8Bi9n9QEJor8GjPbe5xRdVKpiPkQUpEZT9jrRAfqk1N0oJvwH8oJ48
cehHYJid1R59puSFoJuCDxzAddE9KBDcszIS01MhDeYKJIEvLGY4wgCD9rtMPuGaQCc9tqgc70bq
YUU+swGW6bgSAwbDaJmtsExcb9a+DPR53a58CBEbWtpqI0KmBhkyWwSWGFe1Ndri+JesBDkg3BLU
PqjmgZGSoxMkwkoG8wXF+DgPz9PAW2upcokqF6Xqg2U41CJ/EWDrghGVuKB5CD04AZMpotUN7tLg
f8Rzv2Hq+Qu4007jKnuM9tagvSr/UfMuVLLRnL8yRTGiYEL3d+Bdy72wgnVAd3vQlMjkSL9FbD6M
ItlG+HShC/0YSdAatOheL5LmUkO0Xust2EiO7NjTlhGQz7gkWdkHNqZP3Ez/HwKDhp/N/gMX+e/X
npl1DxxfONSI0uPahRgDgep9ezy/hPEsTCZscGwrozemEs2CNDEQ8vByn5qVi+Yr7n8eBEyPVjwl
ZRe/Lfx43Iyh5nmg1kYxm60o1g8D0m6UEI4hoUZgis/waE0KqKDQU06jVJNO11AjKgdQhFGcsqdi
7D3CZBd0tVoTu08hCV2KlSfKAhpo0Y33RyTNH3sy0B7teTfhxlUUTE3DSH+ceHaAXmURQIn5hVLj
8iSIk1qU1kGyxGF2bydveYsxSp1xsD2IRmJybS+uVVQUYBGiHffPAwSkukUSoGHxYlU8R38fi5gI
RnBj5h9/k780zVFYU5ByNIRBw8rFajsHsh5BP6xitcr/YoPkFqghOoDO/24g7eV6HYa+ncb7xASe
lQ071c7eweGl24FkrxhHS7xYuhrpoYck+XU+uwC641iWbvEdklxqiSsu3D6UpKL7xn2+LR3C+7Df
6dGEkXi0aeJtik/Ab3r0Px+/vGvamBInQ4rkuK+BZq7JUlEaQTZ5twemrT3u8/cODyetsGDDiwvf
Azpeo5GBzBiCh7zWmplNGiXcuR471cCfSn3tnrRIV8mzYI3wle7nkF3xaPnHr4LUP/Jk73rWr86j
x7yVN+fdBbsESpbCQx3uIyw/HsKDCY5WETcQBLtNCtRi+8TWCmswa5F1TUDhP27tMsEqCTVWQEg6
mHOvEzWypq7nuyT3078g6vfi94EgWaiQdGTzkapS5jBGWiazKP7s9BwA7c8+CO1/p8OyoEs+O47J
Jz4hO1putgEwgn7slDvtqUPBfXsPHBEoaWlqxhWtLlHTaGTtuI4JzH63RNIQtGsQdOuqHLlKozCV
Kh1ItapbcmGDmD3x6tg3m+ri4cWqiQQSejhYJ8Dl7rmBXg206VwS9REqWVVENADuD7msfRCTpD54
eayq2Fq9whBdDfYUKhu6P5OKGKggq/SB/QEqZQJO4kwEyABDsyfdJ6bxzkNRwTTesJZbItWTa+hz
xAi6s1BFL3GVhPoyyxVDL+2/rZBnjV6khleSfz5rGPesp6C3NPWJ4oUgJFuY4yq8z+Gvs6kF6srV
0kXOiFEa4ScTWqE4t4FrF5tbQ9d4C5SNpaKk6lmwSvXZRdDyB4m0jEswkB2Ofk2hVe8cDfeQuqx6
X5ibC2kyXJXwkvwYREd8J1pNDGLJlu5TVGax0ku7XSYQ1dxf2JBcfZH+yrDLs53Lpo6djNvfqEL/
kQRJKUjNUj2mo30R5pReJmWQpcu8oGIgSmOv46DDkkSjK4MZRn0yt68JOIv7aE8pxq18x9X6gOrh
rClTYvfRdvo8QpDsuckzDNYRcCj0NZLKHqSeE9kJ9YsXDR8M6JBuSgYZwUlr4PeCS++kU5DCMH8W
ZfcKoZxY26D3gxiL/wyRJuhHKMUXGsdapGIrCAdm8Otq6AjcUQgdbyPGss16n8/LehAdFhPgH+/t
ofTjW1iG26drjLdGUmym79p7XAO2iwPQptxOcprT9rjWj6QQ9eVZKapFb24b/JQodmBzSUqb9IIf
OdZz+HG6AmLTa+LwS699bChrXgA7Pj5vODo6N3WmFdGz+nlRYynoD5QUAv/mcwuqKeAGaQv3ToOf
cdiUOd1YppeXsnyvNDmhrDFQxyzHjSWskvGmT/rRS5Ad8QeOySxlD/2AgrybmXjiS0fioFAu4Fhb
6k8KO6pqYQtjm1d/3QMtOL2YWcmfEU7MG71LQ9D/HMXQyA1wBk7FjmUyGzTr9j9EkiGnsnZYQga4
FPoPwNAyo8kEjnFQC8gPbgBOiY5G8AZtCaAqxb47NFtsKY+NYqzhmkRalY2SNXIP4MZvOKNTJhM0
dXr3ajf1gPKRxL0q1pdo9EQxqdvPnMdyyzdFOphzJ4fAy597IAsJZ7nuzk5IBvV44LD6dPoFzw56
VIvezQtClgzTJDPPCH5XjTaGiz8oYLCQ+RaBAFaAapSEKAO7HmTDjOYWnENowHfvgRAgl+FVvEOi
2mR1onMfmT5y62RfX1enUV3DJ4qQzenaviscBvLpFH3uvYpXqeKG8GKiiKGRrEU/onrDqHu9wCIf
5iBEomOkaDGzaqaoyTKxHQzNDNapxaK1rApfgVd40n4aHq10QnrrbET/tVkVMB0pP7AgG2O1/7hL
HD1OFtcwQ6dH3PyB9b1M22YMhFck6aweyYvYsU+mRbOz8B/97AbvyEq6i9nYIZRbJRrAMKN28qdE
OWoFSygVYPfT5MYhfvzevvoLVoOPU/sVcfa4+5oYxuAIVDOktMZ8YmazDcjKq/2HMtkKcwRSVU/F
vq5XNSEr5uyTfPKuS9elzinVWvbvYFHIsHraK81s/Qr/CpWFErKQZljP11bUPH2FudyRcVvAwy2Y
aiVJNSJEC/vsGLXqTfyhL7M6jphL1qwbfajQeENDnbgfS5tm5nZBBEh9w+5jY7/A/zVsNHVM1zpf
TIjxEXbKd/HpRUNqyrrP9Aq9B9srTTXvMD9gW+BdhaAoB93QIO4oh8Wo9IBWMhSAelEUWHnCDfcQ
9WzV4yrSMlmqJmCOzfpF84pGzdjeFf0GgTsGthDoghNy2nJ5kLf3z7XFsOLIh0KfrLhL58Dzlr0x
aWE1UCwq3vK39vMXjlZ7LxBszUh/Hzq2gPjmsDICB0jAgJGUvgBLRL7R12Z/fz6uicKlJhPlL142
L58fgGiQHMEuHId2c5Lm4YLbvNduPYYN/RT36c6HYNJRlSsZuZtIbI0+JhxwFwiyrOfoTMONO3rt
tHNYx56yNm9ZKUDVvn9uRyr+uwbfGNZMiMVosUPJ2YgppnwoBn3eyqtYvIPOmQBDONnPuBl+29FA
P2UU5TxlX+5YDm4+mhQeeCX6u4eEZy++D012qD4HevZBpE7lBDAd5CKiIIBo1Tisuh3lPxzSMjSW
9vPBds2xenn1q3MkA7BUzzpAbp8ovfgINvRJ7cKQfDt5GgpQypFydF7QovxRAkdtYPkACelweleg
K88ZTI7Quf8vzfA8L6aHe+51qjvo/rZqdOC9qTMQlgryabGOTKErFQtxPsZwMkAm2KkN8iR0H/YB
mYjGtthf9acAXYtxPw+hsaxxQzXUWuWzwAJN8c6R/MPLK3Y+gY97jeyPl1P+YhfUNSOQWJHVKg4g
eQJG8oX3pX8vvgXCkUWJXcHXmEAScnfiY7pNTYAr4285UW3hjmL65kHTuYueqkGYaKuCLFeAvDs2
FRQqXccnWpVgdjuOySJDlQsWN0bJh8VpqTiWEFmR4DfDDRnfBCphW/WdpU0CtRAOk3tXgQm2kkwL
Eh8e5dL7IRsfTKOfYyNnW0TfGjCrwsBSmUN1M9K5oQqaacFJfA0E5mKW1BSvlrD+RE3HhvDUKKDU
e1Yb8EAAjdOmOumpwE4UEuwhvCTQGnlcimzqGF4oSANnO6CoWqcUr1Pfgbtk6oI3Peckymst6dtT
APSQ3UtKD6gCYVPlKEEAFGFOiGOAOlFgKrC9eLKQTHxfoYjKOJPgg5u00JPOz8y9tLQ+RBCSgJNh
VR+rUrm72v8gsHLvQJsP6l0zWc5ZY9q76GImwSUKD+22l7/6SfD5bX+LLdwaRBDHULtX0emxGo/w
KAbFfgbNOwoMCotlqenR90Tks/z/2dahhFLJNO/L6AhvirYzhfQkVt/rPxWjRWaLw3Anf5isKS3L
UwJsIrvAgD6ZbiuYoWUo6SjmBwt5lV4lUJ8s/H7FmrxuzwRqTMc1EKP8fpZJ0kvRv7Fzr/MTP2rI
5SNZ9hSwhf8i88RyIcG9EKC1QUxj0wRmCl1qu2Js1rtWSq3BWyenqzGwPe6wULqvG1cFWuYeh55s
gsX/ArQX6Yq8hogkW6yMqEMj2drQasFIBTvx+6a67to6nWVbWWr5mYBkDBMRmuuwCiOPCD5TPAvU
RyufESZrwzi1DO/lpzmP7kK3kbvo2igu1oIaht+Omqpq1XTSpP8rJlQ/YV2wfXuKX/AIU7kHF9D9
6bxVjrdLdCnkZlxvK/dsB6nYuyYtiZcwpTT9tv+DCMUjl40onkQRWpYwTISNirLTDdFuYf+BdmGd
DL7D1bH++y2f3UEecQgesD5DIsrY8/bF9PRpVJoGQ0QSjWxNB3DhuCMoA2Qtkromu3GGv0m1d0jm
VSGlqW9RTmWCThcz+6jpjtSjbJw8IcUWIRb2X63xP0mfUOdXlZ+NYiOmeDQD0wj9NDUWPr60eud1
ezS18AuUWdD5N+vTD0MQQ/ZPVIhipj3m7rlrNPBKc6eB5DShdG8LOD9d7psV+4x6Rq9EVJwuvWum
SRXtUCC4TfuQznf9la6MvKLhw4mZb2itog2nrN2bwkStpvICWUWz6qrDhRB84+I5guW83WxYaR7H
Tflu34/oCVgPds1Z40lUZ9Wr2Xy1dAfao1DSAavRtxY5fvWCpgPGgv3wiL8CX4vjDoFN0+SW/yWk
0C/uUlXdfzDJZVKJFaPysfXzhLMxC6k2x0yhgI34hhL8WOAdOM9GiaHMAmfrACoTK65B8GrFY7FG
p+L1qQqId8u4ZNtPjkax8uLd/QpNM01tAB0jXJiP47z84YcNPY7wkDY03swvYBYmmPadRyyuEHDA
R5xysnIQyx+lhpirEjT+S97TPCCYySBIU9DiLJQqacFVzI7YNfX+2mAXtwRxlMysa6DXunrCz8V4
84VWTW9GQ6F/HhiXJvb+TtQ+eR5G22trXgk6yV+T2qwISFH9pfw/EbP5Qzofc5e9b6+cRdSayRVY
Zg1JYpKDvMCQsc6khSx2vI2t+u9/axpHEoKrtRRE4w/jGmGxPs79gizzDlbZTyIhHAX2O5lTUcFv
OyJQvISmipak+kFKTnY45DGuSIT9dofSTAgnqHY458f5gJUfs4X/htnHuqNjTNqLTRKEx3kZH0CA
GpCNpL7JyRQnehcpslHn1OP0uqxXHBv/hiHE3iqU95ps6ALZOD6BDbAyB1y9FdpCRmzD4m/ubJy+
di7FdgLBT9J5ovcAjLlfkuNShuTfrZKPs6JtSLsDXKwkJODmxAVgozy15c8uriff/YgWL+QH74PB
/S8kyqxwkgDmgUty+tO32hmFfcwiqdfPQciE+Tvh75LaE7i6PERgwVZmfrQGllvpUlcLHLmUx2+1
Ni8pBeRVMZPamZncMcpqJmQXtvepxM2GBFT2jIYInfm4dWKccBN7rJmJ0rKMHWDkMUB/2cyL+Y/Z
x2MegeMrJGgynl+kSZNZmFsJpcMn4feg1gU2N08Hd4ve/w7ID1WIBv8c4ew2vPSErAErKdLtqVM5
Pis2DG6uG1tyYzrFmvX6E1kftJdPVQyIdN3aFFJw+0sVkM1mO+mMcuu2+ztgA2sPMK/+x/e+pbub
xR3ZMtA78mrMWFEMHJSUUBvVOnuxGahFSQR9KixbehDDkX2iyRtEcKSTQYEcjg48S6e353XxuS7s
eRJesVtKJDJEAlpv/RIjkeEOQlc574G/2HVadhgdZleEOyrdpiriwiB8hBx4Baeg5RzM4tn9ElkU
vF+7IBRnh4MUNqNhS2dgjlpBuMeTKoSK/UC05ThePgwIuGZwCM7t6WCgjSLqoQZ68S0atfL/7vi7
bESb1iPE6U7hvz9xQxkUmUQLLIFQzpmMEdwDp1v0fG5TdMHIZxzRJ/Dcju2jwGuQXpwXkc86cZIf
sH/t8w313GtHajj7XT7jeFjUXwufSRq56YqSatb+XTNmPcdoP6xFUirRxF7ua+8xhSv8wSdRoK+Y
HR2uvqmcr/A6zIGg4k4jaRm5yYVUU6m0Lzl1nKyGO3aTTgUKWtzA1B7fhN1NbWeIucyifwjiR6OH
crwgZ1WW4zt/kzuaMLf1FYGmEV6sppFtQs9oiKFzR9EhBtfUnZx8wimoYhIQ2xQ/dHtfpEIZe4vq
f9zhB6tCJQItVGLLBLsSIkWZX+HbDVF07uPxReIZtQdekFa5n8BLEvBkZJl5T0hsPHwTXomEUGPJ
HJApKP6lgrPK9Xx8zeRIvuauYWQsT/ngQjFik4NyjW6s5XzfKKbykC5+zQvsQS8FyJrMJE3QDDRx
4smCWEIzG9OjZlEDH2XEK0P5n19zrzit6zh5ZESCQc35BdSGlBky+S/I9tFfZFLz9Ku7rlqJ/1zb
b9ubaXyAhXtfZmB44h5saba9oqdtDUMtB4j4lx/zT/O1U/hL0BBR+jJknj0h/Znd3vH0zaYGeHTD
zZW926fPouRKI9xzOud2CHd4M+fSf12vUHa4jB3j4Mi3lWM7XXC2baSiyOvai3SRJ1LMUjg0BXmw
mYlq+iShIXWV+CMRIdOqrfB/nLMQYsY+XrrZ+gud1hiN+IxOECIqyH1vPqLUohPP6iZzBWYANZNJ
NHjz8y18NjPvKc7NIFgkQRGQa5AUTnmws2UBoOvxebWCy/tTOZbwWWkOFko1ToXiNJ4PpJQQR1tp
3YLZqD1dniZbw1WQgR0wrgrusFxiyR9NDU+fV9Dc1DImusgqL8sH1eBTwAMH/WA7nE61wP4rj5YB
4xKgDMapKr6C40fPFkITwaBkRcJ4BNABH62BXXgxCnm4ujTMkyXDTTaQ+MIh5xV2vaCupqRrbOqv
eSEM8vmRCXFiu8+tNn1Mq8W5/vfVhto8ZjGCCzj0VqFQU8ZBB/yL5g4ZRfnVmiTNYVNd685jQiyD
5Vcu0ZxA+uoO4U0LIJGrXD86V/ozEvFmZaTLwYNOACqReveWcNyehBkmgt8+zcZmu4pQNWIQDOwe
zEQUo+IXTd0t9SN8NI/XIMiKr9X+jz8yVQpjtFoOzxCqh3zkOQZwThPCjCFuY1omPYCch9/+TuL+
CyG/5sWi9fK0reLNRVUp/mW28AD+ubBy19YgL9cQw6hvMaBsA+x2pfDtNywOGOBVtLVfWeKiQ5cH
J8huvCs9mrmYfbAhMkKvxf3tj9CkBhKZrJT/+GNG3bFI7OR9lT6r4a79GsU4Cx4k760sTxGUHCP2
7PijCxulQJAD/uTgGQMB3udIe39gfn4/7oX3KBaOocRuHgVAgWxbATe2LverO67J85Km1++y+8m2
RfN0GJeOtCjABkOioqBD3eAMwLcJt+4E8a1jqZy/lvny6LNboOIECOVPxA==
`protect end_protected
