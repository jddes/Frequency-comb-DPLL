`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AJIbPqECCn0bmGxsdLM1onvC/TqHTSF4JPBKyazi5Tiz71narbYuqZZedsopfypdXeYxbli+96IT
XHSEEyyuzg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iD9ZnLfSLtR6+EZLSkLC4pXQnP0vlxOwOdTekH8QqSan4Nom4qzgcGtE98iVMOsWGSG5K+3+l+Cu
BY1dkz3XT+4bRbL5bYAC3Xw6P51gUQElvpiD5x1e9SNbIzS23CTsnhiB6p3aCKPO2dx3B8aZM2R/
Tzc1RTZ4OpZnk1XY3Pc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qu16ZYk4cBn1ipd/oKDaC6S8krPdgXVhiEop35Thfh/zhalGQDF+nuARPQZqgw7u+5QoFfI7dpcr
AkVAZYWRSkMs3lyzqEcoAIIKlQKu3aZhymQKA/d6QFfziL0zl2Ja0P2svGqnNMiGE6YPLI2bRZfz
Zv/ioc6xFU19QRz6aYGHGrhGs/dnqE7SxLsTRsPobdWcGOuVfcf42EYge98WZU9uhJmnteo4vPHV
TriiOiGSGMqncBUc4Nf+aeOKvgLQrhPr6CdvNgMTk/mCiYxaD8ZF7PNX+FJGNOFV3MaJDvVHE9N5
W5WiXerdLXuo1gu5LCC+CR0tEdgbGOQR8u0vjA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l1t1J2vI/xDoq6DIdl9ADGp/xZaPVTscczRj7qsLZA3HO4sT7Ie9O/b4MNPZKAv0c/+T+wy1L/zy
warUibv0zs+RkCTKGKXmH4WUoV5mTe5TUlGjIGvgR0mCpOK88zVM+j2t8SEQUrTYbn6Y4GkxSTQf
II8bXNd1XSojdLfp/vg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Vn1kzbTLA2ZSG1wKdTzr9cGYMzXtCSgS3lqKY1Xi+f07Qbwmil7YwaGQbJwQledUmX91HaWuwWrC
tePZb6hb1vxz0hby/7Aroin0LJFc3RfdTX0VIcie28wTpEJjcfsoHBpzopqtFMBm819GoS1xag78
bgwmqzX4vIEtTdFxocV8X6XsFrpPS3CWRBEVs9l6gIqj+0PHp8+Z3sdPn+16DvFnlhD265d4EIOs
f/vokG+mWlHb3TGFVFFlRgqHqXZFyHs9fvnWrID3/U1+0z2EIsVSPXxluah05QLdFF/CXiPAukqY
HANVxghFIfGT1fZ3DVSRiQ1Om0bJThlCcPaWTw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AZuc9OHyYugQnrL5ARLUTn+MoogZNR+towD1VEaN8pgKgH+NbVHBe7L6EL3mFcprbbAkivhAxr92
jAQpBGLqSGxuWErL4Ozcc6OsmJaHfc2SOlSgWtVflZY+eS+kILpe1EwqWM5FHQl6BLinutHueoq5
idnkkQuCiUoDbV+LrB8FieCqKcPJq/CTMfQTFdEox0sFw2N46GuZ0Z0zdHphXeSGHgSVq5r4L9WM
NRV3hevP/69Lz9uc/YB0dDS1w+/HBK/WTxgiOzqGI1wm+zNwRpSQypY5oC3wR5jGSKAmLDOu8EjU
FJAFBILvzYo0NMGI3avYb9fRd2GRAiYO3mkXow==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5872)
`protect data_block
/QzHe+sQSaqBa5gwFdpGGfs1q7YF1QTFviFwvSowtJ/pgG8GPo1bWLfBOVWUkHHRkCISRYRa8tjR
CEAOLsnf/z8b2RrK+5So4I0IeOi6bso7e6yL6+ojfnbXatN7U0yYjPfdnVqF9omklMr43ZGreSuN
cnHrXNFQUGgKeCXJppSCCHM7M9OE80MRO8W5nPYz71AGdlH6jgkr5J2rA5dolBQH+i5M2ZbuLb5x
tn/1O+nxrGAMdfHfgPxVxscuiIBkPawDQHD6/lafUBYlKvIRJkk7tVTsYMFjKxWF/LCoJ/KJ/nYm
C8GXE7w6O0OJN2ffatIynJyfiSCwnhukp+ReLnYmcgU8r7dUzu3G5tGW+KQdpC2U5xM241uR0Qit
1LUPIQ+aNUzigHcaBl5bXqB+0xrjf+aUtDjijJ8BmJssQfR4E+uyMZKH8pd2+f+48uZ7rVFLs/Gm
IgZXoHT/GwpXE+lImookgOGAw7qMahuK3zQqrbkrcMeZ76qHfcZjjCOIEhHOaAPnaDHfRgC1Z5D5
qdpZJQlUJIPuAlhNrqVaA+eJjG+XsfIBZbXGSTdmt5OqM3KUFnqb1p6cUEKal89UbYHlQjorz43f
kxus31slpxSoxUNHtslEZz/K5w5e/2Q9M0rXHm5CM2T/2Y4VYyzIEymknVWghrracAaxkmVn1RvW
qWwR7RWlWNp9ZVQTuGbg/kMHehLxpEpoLNeh2VeTXii1SjRm1epV7500CpR88ydqAlhAHarL/HE4
mTKVgeXp51Gqog7wJpVBany2NNcV3iPJqsUDzwEEOGPCTaAKMWgYG1xKxM4D9d4tOII7VAFfpxJG
0PmjseNdMZNonCkMHcSmuS85BUxuh8ig9sdNJxYhLm5OarH8oAYoICGOBg6R6T+ZW0CLys8rjJfX
BEmYEzhJ62/d4gKpk4FkzydUMUU5X+sQzSOQ1kH2WmvuVU48VlE8VQt2ck7rg4lmRsisG651KHCX
Jo5vQP/nVyT3yO2ObbZy2KU5CdeY5msS7AJYSgRShb8pWq/enU7efKRc8XtOyO6a4xSG0kDN2wG7
YNeIbenSVBtKRzctXSnQVSyGZkZr8LYl1wBvjGBeqB1hqOpHYXQNR5Z7kiXdtQv9pCVjWN04r8gq
WSUaxkcKtLKRYkcOZ5IHsyqswB2tjkJnBEDtzck/ZrE7ACTvaN07AwUvUHqyJ4yFSbqNxobqu+p8
zJ4mUC5eqLgQu8AGJg0U32n4i4M7XYEAH8l8oshyXkrCppT9Tipkc2bbiC0Az9UBWYCIkbFbL2su
F5ntqh5mmR61bRYONbxIrtx4U/fpb1KT5ZI98H77d8GTCjgJszJu30Q/LcvnIyfM3BhE4QZnJrTb
F/RI83hOOdztFwbqBJhSTl9gQoRXeUz6J721Y7+S12G79MaGsEe47jhdP53HVgwQ6mRZQyMkSB7v
V/FDT3kJSK6nLtG5nrkJGzUHD25clSN+fThcmyL7n2L5lcl4oFHeCjGreYjdWgpz2cx54KEQWObV
uFYjpeKvJKlaTVdZx1P+iic+KezkQ0JNWLIFJ7kbhWOQo1PPeunVjxAq3Rpcs0j+Gnp2ivKPL7yO
t63JkprY257wnVNd8XWJnVmrlhngAO2c9a9wWVKw9TB0l9oBsINpfyOFmcXLEPxDP+pAPIjrUiab
v7jn8v8ySzSq6ALrrVfD8GylTz9KSfbpgblvMAuMlK7M1ihZX2H5Gi25UzrgbJt6iuJSjEpbGfVb
thDKRjBtvskjEfKkKAmUQFpaiH7dHT87lccy0ULAHEePKpiaJsjmlzy6Eh8Kvjn/AO/FLJnNRBuE
hoqN6kYPQu/QbYslEAZAVCqdGhZlOPAORzTUCYD4aU9HBHyh0GkUZCpvPWN8x7NoqJHjm/P006ed
jKNii8sQPDnFlYD5585K7PrtFdO3UBzaWYIvOr3I8MJAO/zvCBi3jxvjY/Q/Rt/Y1r76cqCKPhkQ
+hYt1Ftmpcofcvfus/lYvOCh2Bt+tDlZITXcWCb6XgGSutqfTwOCXio9WwrUB7kOA0y5ug2XNAqY
as52+m93y/yPh1UxXSZulS1hY+hhw6DUKT/iyaVPqhTklvAsD3T+ATFxE7BQgGAAj2C4LF9/EN5U
+CqC/i1GTlKyzmhsv7pNNWaCn7O4h9NbL4WMJdtoeICi8ZwjpgWNqFG4euLfCeOf7F5x8LsXg1cK
ngNVY5dseDr69ITQRMtmTXxEgcgVCVRnyqPwQ4TU6c4tA1g+/D+Ay9xbYJJkhCeTtkJtyppPGXBN
8D+No4T48tC6u5eLEvd3X3NQt+Pw1aD9/phQ7EV9+ZIxcsMyXtfdPSq0Qt0ny8TrOHYBBReRGajP
e5dD9ZVjM7w91JFDkckCgh8w5jzn8KOoGSCoqaekvYA/1b2kH8d7SIHsTGEt9ahwJzf4+ZGPL3P/
veoz7P1ysTY0P/rcjKHkJbHJ9RfsALF0szoTDZDhe5afyjEofUrRmmvRGXaeClnuqEF6xCQqku4E
ZBwkmREq+qLyDldxFnJPRyFk+VagvgAR+F5c3iyPnY7Shl2YgsEh4iKr4QlehPjpbGiSY9XIDBf3
yZhSKexGSS7EPrfLNBOyOMZE1Gv9I53jWwA4sPQFU1zDsiVwk1o4P77TogwQf2MEPwQVtURWLp1s
QgxQdQlx0gQiAiSIcF0aETf8sIeJ7PEQmpcBHsP0ZeWPtR5FiCr9+fM2K9nKB5ob8OCJnzEnK/sV
HZo8GvdPQqySq3CImEpaMFwhSjoR9RNKoBBj4Xy/M1PUL9zFS/CaHR25ocvMYckgynQUWO4d9L6X
1etTGzHxPf+wMyiut3FohAJ30ef0kTDISGneOvE+obT6aDPZzXrXwvH+4POOrKdfDbQ1VJBss0M1
HXSBk+4zcXt5WtrwdGvooQyKTAhTwivyCAE3g/uleOl7MUwPk97cYdwMrMiDPn7ryZxQAEdQpSFK
+UOBYCk0kLaJ0WClholuoI4imNGgrnqbnSF+PjitTq2zDVKzQBUDHo4dHKEgnPFNFDT182GjXwCW
t44I0KYWiDIOhEBmK/zeGSG1w0Ut+lKh7nBAu5zm1Jh8FdM550lJ8GdgWbVcbzBWCef6teEW/p9B
e9rYqLqVD2KJYa8WbUhd12dQTM3WxdH7maeJqKnm77NU/RYOuiZc1BwwCn3zB6FXFYSjFmSnqg99
s6eeLktO8OIWMsTwLk648rwjtFFt23kIxdK3Ibc0pxkpNRbHf8gUYyOJGL8ikH4tOIhsCFajiWHJ
vCtpRUR5fATd7UB54nPrnRBKOjKCvEzJznOYdWhltp7dI9VWgQAzeimkfOT3S2QkMPOsYTTLZTX5
Pp+Wj5sATZexVS4o6GEsLniqcvp3U29ogBqpHsrg9o1VJT2rtBgUnEA3I/u1I5D1V+f/r+mnmdRh
bXRUjaQ3dINPi2LzZ9eBchWHytYtwWfXOg183oILSpenj5FXBA2c9LYMZDaTolf0lI/M2X/4AJwW
ku+4g3HSwDn3bMoEHTcy1avO2jgeqWR5LsyRh5M0R+psSSMDLNvDr9m/Pfpem9kA2NjXZfWrKYBF
iC1OTpkkizU2wsx2kd+PFcF2WCbK5oQK9gl7gJxFyzg+MQUq7nEtvrro8eF5m/v1DunjAevFwkDc
fjpI8/lRI8NFqxyF5SxL0ko4X8yJDCRmymKwmrvGP9vueoFFJQgiHoYap1MKQIIbRiJrEpzyPi3l
HTkeiqsnZms0Yy8ewc7orDqJgBmJyuZXD/p6GYdAyLJma9xGFxh9FtTvo8gXBE7F2Whq5jbvye4g
2olzRWtCAiNyjsdr5GqKNlf0um3lOleQUIMmVdxBXRv9D6FnNMEpiMpceq0EnlfDwP9yWL14ed6q
/pg7Si0Zc2SWeKpPziRsOXopZIqjJj3sISCvw+dtxOCElX7nqR4GKhhHCPDP0DGkloqDJsgsqQm1
xZmi9SOrsnD3WaaCNH0PlS/DxOmtZjurUtDhINVJLePLjJXgdXHuiEzl+ibC8yVxw0g16OOoFdoJ
JVV8XXZ4BubYtsoAYCZgMXzkTkSyYlgEUbnpcnyVbRcPZJudT2USOI8CQmYp3746vyM14fp4AARz
707BjYnUwbx3Bv00WwdLdgUM/+ol0LrPKJg+rUMA7iqWlL2gX8uztqkqhOaX8hTKcPP2eUSJt9tO
+9nG8siNCf6iLXob1tJcjbaAeFoW0dcCHZ7QQrQ7XaPKnvASAqevHsbyCe6xEYgJGCIIs6+CpndU
yRPwGsv9rX0VbQrQkMWiZnVYCvA5kTH7115Mk6v/ecgFng46OGnhiurZAwklPAPrJxhbIC5Ni4Ja
Lkgm216ALlrdzMgmy1tt9F2j73lD0jydjQ9M/6UgGxeXMZcZKztom5Emmd/mhgJ/iY29bf3YegYs
ZyuaZGhNqvcl0zTSnd7xenxP8UJnEZqfmISs5mG4nJsOx0W6qGEZEwbKxzE3mK1jfpi2uJysFhtL
CS7T0XAxUqVD56XITwLd/CiWlr+dhqTd8mVrQ0xkbf2bHPjAixkSwlPH9qBcF5KE7x0NC73rllLd
uoAulxm2A0P+TqBEJQSOqpqf5WDd57rEfiiP4CsuEcIgb2yameMAAYYIe6bB7xJ1GZVenGO8s5uF
HCnItFwJDDdg6xKjwkcQXJBzC3z8JiFquaVnKz4DTB3qBzN5uItxa0swaWleFK02LhEQtl8W2Sdz
pqgb8CgcafeWS/faQZAG71GeI3NE/n7+NVAtZ1FX+w6Q0v0Q0X/MyXdd2lI0Tvf50JoV0ALLI6eO
RDdPAz4RhZ13zIatxJlHLrUDJFi7NSd/NX+wk/RRAIAp6B6SWdB5fCwVoPGhUWBrf48dqLKRazy9
9JasCFDn+hp9TV5F9yfKicNkAwX8x2yjKEKwrqodrmQZNhXUIMUMzyRmEcK6uGEj5A1uyQtldTUU
y4PpRoxOdNcZdI0B5O2FhwB5H3LbhPRf0ZrNuZQtewYL+c0H6sPUBm79zl08CNl/jTguaUg+DpRk
KQDdiP6W39Pa7sxN1OU9gFLFKDAOTLpmdgY2bDFYdbO/0TcusYjL5Zkj8/CGcslPn4pePK3YRhBm
Mg1JK2rM2xHAQfQeYvZShyq7KRYY44JYnE2UAiTCdXuqIGFRrMakQdcG1sCIBZ6NLdX1ad3KzYDG
/ySgP965uqXqsi5VDPxUECRXZRE0WHSaimuSztuJI/xLnt8AwDp0iUaawszKz2GnNRU92iRHcYoE
ywd/k0m+JoltfQYxTVbdwOP/Y6mU8TOFhlLZOKvls2ToGybQ/2ezGbAniiliHa2nkLtk4IxjfvPx
Uc2hbdFalQW121DP9r+Yw6Uy2rMFGXHFdIGESPniX7v2qjCKNKQy+qRkF7Q+cv4wzzo2ZBj4g1tL
BWKsFY8w8F3OW4yHecn6EDmlYf2Sy1MpDNJwpZD56YJH9o52r2IUJUnr5I96pAnh1WAGQbFDMX8R
HCXRI7wq5oJ4hMVh7JBj8jcICtFRrWC2TKtyWD2fBNFb8TW8+YDSqIKkeFjctffgSx439NrFIcww
3T+rje8turjFg1VH6mFQNVCbgCQOYeMr53WDtMpsBfvl4kxaANMS0E2XsQ2AuxrHpfnzxaScfUHy
4TDXCxenh+8WK1snhHRDhcOm+gP5aEujS+K+QAHj8WP9sN4DwDhZ0FGPniTQLxmo14tVg8CByU4r
gZJibyFEWeSeNWC1ik2qljdU0+WNF0LZM/xNso+XKPncu/Z9uQFl5Yn/+0RaNEBRy/b+2Tiwfw8g
U6zu9Bxhls+EeolcaGD1RB/424nvyzpYRctLNEWquVXoQwyNQWXfW/i9WB9yXL5FcLIVkM4qLqa6
Ug6n3RAZ7bS/ect4to/qUDvOp0ZznWhEzF154+bHaxFxSDWgz0KJuim+ytdEwd7vidKzWdftKVjB
aj+2ORdSLMOfgCA+N3xavuUCnvD4W/a9ZeEx4zL2e7I6XBBkLHBozvVJrXrSaeNleyg+zTNCV029
M/thKy7gDMDm2SFlJuLBmfh+/Jk/Wybp0cI97/tCZAH350VFpae5egbxBc9xhOZXoBqpIVtgAS6g
E55XTJOo9TIL6+sPo0Lp8oy84tfEADNSW5XsGQagQOPHgLu0dOBXYkr5MOew287v3F0yxntsh+U3
ZzWFiWbjou3Hg2hCUrDfts9T+9QFUZy5HsyVdHtnd30GjPB7T/Vl4uVL82J42c/6hpNRnRu9CScz
8j0+x3mKEzs4I2eJaMHiRNfUveN5F7lWy5z8H8o7zobCDMsI7+9iTENTKkniuLUsuPKoONG+gx78
LZEF17uDkIoGVpHmj3KjLwZFrld9DrFJIoVXAU1IXJafJjRK4n1wRrLrN7uUgCEwKYaBw36VJoYJ
1Dct0rkAEI+JWfeTi67uuS4jIqLGkzQ3gfhXxEU47SQmLapf4wdf5OSd+gJVuW2HK9izBj4oOrKf
PdXbcJlyF3TQ9ch/dkVVdtNE6ep0BozMEjWQoF9aHD+Nex96xGdNDSUbycptx8FmKE5dawGQKh4q
mB0D9mocBaZFiIkwEGz+5uLk1lMx2k05DoDEC8Fi2tqOHnniF6t5pSa84bDBeIrRO0iownmAC/vM
BsLXijfIIHfbUn+o7e+UKxTUhphVhv5tpRvplL8YmTxOmfygSQaWIIhi3DeyuI5gY1mOemyLV/SS
foo9uS4ZvQUxW+PN62pF6z5xGrUrzqAZ4J/rq+WJTR97d/mRMO9AzuivyiVwynXSB07HT37F2/D8
J6awILrnSoet8n4aB8vHHvOPDrAHEq/qrrqKM2HgCRWNSXgMLfDddrhIBGiUiQmf6mm1ZumJ7pPS
jSy1uE3kEcxvAMiF1G1n/VfDDptVqekAZTHTlU9VkGH8/444j5S5FkYHinB1+9MSN+ueflNWCf/G
DVt5iDfJ7pPhluMzmg7VlHvHJQ7GyGVal2QqRssxZXb/aN6A5AcEZQttgLBHIOYQ9HHo3X6osLK0
CS9QMiaAzpJ8RawWXTvgNOR7cAuHkxHMPStUnlJHIk97QqdiQKxOzJ9vLz50I2/4c0KKzP/XBzLA
Wu5/PeKZp8WA/mkurTkd4y6ggm3iXqeyNoxoaX0yBOieBz4xDdUHD24btVoLEFnPW3CbnsGxIYRZ
2/H7cNXOx2AuHe8Aay5+ke2S+GeJpCUlL9sbuyj3ucdlOxchtgi8yL+DPaR7pABWc0op80dYxW3d
y/RzYbuLoAW3++1cgcje+vpYSLPep+NU1Qvc8oF2cw1niS89KZRl9Hv2AZsBbRdSxtyoW+7SS0gY
/j202BoJQ9C4PLRyB/IjdyhSqyS3ufFadqI8NI5lB9eD0WT+tJOhf7r074frE3Q1YT/nDwAVyubI
9OmwYz37NxNH+qb4yor4fJzAFVuVonkT21n1VlkzYxZKHmVt8aoxIXV3pvCEHPNCDMrNzoUxR98V
y5fiVXa1D/ho4I1BL/0X1jFhrIWGEPs+iuTi8CmhYZGSt6w1Wize0LkE0LvRUYvdm/snUU13GWx/
RGhUuhMLLex6S25UMuLoiwHwG0eH8myicWj0691ZoCxp/xuDwvMRgz26+RB2vXCAJcgpPd9fxoD7
uaXqS7i1d6u9Lm2RtMOIMLoN+swe7UiWiTKzTzKII2ZpmzXg6WzPTBveqr9AeBvHR4GTcVPIWIAa
gZ6AhoxbiadFunRR1Gv/t/IACXEfCgFzadV5WWNC0mg5yHQCzGcrSE5tS/Q2cTMiUacRMxSKL9t/
iUqUKLSfIytwWkwKcMtJXNhwe70A1HpnKyDbH25Bby6kSBqikZ1aN+Pt2l9NltmjU+O+cZFGfzS5
bA==
`protect end_protected
